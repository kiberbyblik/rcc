`ifndef RESET_AGENT_IF
`define RESET_AGENT_IF

interface rst_agent_if();

  logic rst_n;
  
endinterface

`endif // !RESET_AGENT_IF