************************************************************************
* auCdl Netlist:
* 
* Library Name:  SINT_mkm18
* Top Cell Name: PLL600V3_m18
* View Name:     schematic
* Netlisted on:  Sep 15 13:13:33 2023
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: SERIAL_LINK_mkm18
* Cell Name:    ENHSP_PLL600V3_m18
* View Name:    cmos_sch
************************************************************************

.SUBCKT ENHSP_PLL600V3_m18 A B NEG POS Z
*.PININFO A:I B:I NEG:I POS:I Z:O
MMP4 Z A net18 POS PHS W=4.40u L=0.18u M=1
MMP5 net18 B POS POS PHS W=4.40u L=0.18u M=1
MMP3 Z net15 POS POS PHS W=2.50u L=0.18u M=1
MMP2 net15 A POS POS PHS W=0.62u L=0.18u M=1
MMP1 net15 B POS POS PHS W=0.62u L=0.18u M=1
MMN3 net3 net15 NEG NEG NHS W=2.12u L=0.18u M=1
MMN5 Z B net3 NEG NHS W=2.12u L=0.18u M=1
MMN4 Z A net3 NEG NHS W=2.12u L=0.18u M=1
MMN1 net12 B NEG NEG NHS W=0.52u L=0.18u M=1
MMN2 net15 A net12 NEG NHS W=0.52u L=0.18u M=1
DD22 B POS DP 1.02e-13
DD24 NEG A DN 1.02e-13
.ENDS

************************************************************************
* Library Name: SERIAL_LINK_mkm18
* Cell Name:    ND2HSP_PLL600V3_m18
* View Name:    cmos_sch
************************************************************************

.SUBCKT ND2HSP_PLL600V3_m18 A B NEG POS Z
*.PININFO A:I B:I NEG:I POS:I Z:O
MMP2 Z B POS POS PHS W=2.50u L=0.18u M=1
MMP1 Z A POS POS PHS W=2.50u L=0.18u M=1
MMN2 net3 B NEG NEG NHS W=1.06u L=0.18u M=1
MMN1 Z A net3 NEG NHS W=1.06u L=0.18u M=1
MM23 net14 B NEG NEG NHS W=1.06u L=0.18u M=1
MM22 Z A net14 NEG NHS W=1.06u L=0.18u M=1
DD38 NEG A DN 1.02e-13
DD30 B POS DP 1.02e-13
.ENDS

************************************************************************
* Library Name: SERIAL_LINK_mkm18
* Cell Name:    NR2HSP_PLL600V3_m18
* View Name:    cmos_sch
************************************************************************

.SUBCKT NR2HSP_PLL600V3_m18 A B NEG POS Z
*.PININFO A:I B:I NEG:I POS:I Z:O
MMN1 Z A NEG NEG NHS W=1.42u L=0.18u M=1
MMN2 Z B NEG NEG NHS W=1.42u L=0.18u M=1
MMP1 Z A net3 POS PHS W=2.20u L=0.18u M=1
MMP2 net3 B POS POS PHS W=2.20u L=0.18u M=1
MM20 net17 B POS POS PHS W=2.20u L=0.18u M=1
MM21 Z A net17 POS PHS W=2.20u L=0.18u M=1
DD32 NEG A DN 1.02e-13
DD31 NEG B DN 1.02e-13
.ENDS

************************************************************************
* Library Name: SERIAL_LINK_mkm18
* Cell Name:    IVHSP_PLL600V3_m18
* View Name:    cmos_sch
************************************************************************

.SUBCKT IVHSP_PLL600V3_m18 A NEG POS Z
*.PININFO A:I NEG:I POS:I Z:O
MMN1 Z A NEG NEG NHS W=1.42u L=0.18u M=1
MMP1 Z A POS POS PHS W=2.50u L=0.18u M=1
DD7 NEG A DN 1.02e-13
.ENDS

************************************************************************
* Library Name: SINT_mkm18
* Cell Name:    scpllinvsl_PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT scpllinvsl_PLL600V3_m18 A F NEG POS
*.PININFO A:I NEG:I POS:I F:O
MM1 F A NEG NEG NHS W=1.04e-6 L=1.14e-6 M=1
MM0 F A POS POS PHS W=1.04e-6 L=1.14e-6 M=1
DD7 NEG A DN 1.02e-13
.ENDS

************************************************************************
* Library Name: SINT_mkm18
* Cell Name:    scpllochk_V2_PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT scpllochk_V2_PLL600V3_m18 FILTER FRIN IBIAS NEG PD POS TM1
*.PININFO FRIN:I IBIAS:I NEG:I PD:I POS:I TM1:I FILTER:B
XI17 net24 net1 NEG POS net44 / ENHSP_PLL600V3_m18
MM7 net34 net34 POS POS PHS W=1e-6 L=4e-6 M=1
MM4 net93 FILTER POS POS PHS W=1.66e-6 L=0.18e-6 M=1
MM9<0> POS net46 POS POS PHS W=1.6e-6 L=2e-6 M=1
MM9<1> POS net46 POS POS PHS W=1.6e-6 L=2e-6 M=1
MM9<2> POS net46 POS POS PHS W=1.6e-6 L=2e-6 M=1
MM9<3> POS net46 POS POS PHS W=1.6e-6 L=2e-6 M=1
MM9<4> POS net46 POS POS PHS W=1.6e-6 L=2e-6 M=1
MM9<5> POS net46 POS POS PHS W=1.6e-6 L=2e-6 M=1
MM9<6> POS net46 POS POS PHS W=1.6e-6 L=2e-6 M=1
MM9<7> POS net46 POS POS PHS W=1.6e-6 L=2e-6 M=1
MM5 FILTER net73 POS POS PHS W=1.66e-6 L=0.18e-6 M=1
MM8 net46 net34 POS POS PHS W=1e-6 L=4e-6 M=1
MM0 IBIAS IBIAS NEG NEG NHS W=1e-6 L=4e-6 M=1
MM3 net46 net44 NEG NEG NHS W=1.66e-6 L=0.18e-6 M=1
MM1 net93 IBIAS NEG NEG NHS W=1e-6 L=1e-6 M=1
MM6 net46 FILTER NEG NEG NHS W=0.52e-6 L=0.18e-6 M=1
MM2 net34 IBIAS NEG NEG NHS W=1e-6 L=4e-6 M=1
MM10<0> NEG net46 NEG NEG NHS W=1.6e-6 L=2e-6 M=1
MM10<1> NEG net46 NEG NEG NHS W=1.6e-6 L=2e-6 M=1
MM10<2> NEG net46 NEG NEG NHS W=1.6e-6 L=2e-6 M=1
MM10<3> NEG net46 NEG NEG NHS W=1.6e-6 L=2e-6 M=1
MM10<4> NEG net46 NEG NEG NHS W=1.6e-6 L=2e-6 M=1
MM10<5> NEG net46 NEG NEG NHS W=1.6e-6 L=2e-6 M=1
MM10<6> NEG net46 NEG NEG NHS W=1.6e-6 L=2e-6 M=1
MM10<7> NEG net46 NEG NEG NHS W=1.6e-6 L=2e-6 M=1
XI13 net93 net66 NEG POS net2 / ND2HSP_PLL600V3_m18
XI16 net36 net46 NEG POS net37 / NR2HSP_PLL600V3_m18
XI12 PD TM1 NEG POS net66 / NR2HSP_PLL600V3_m18
XI15 net2 net37 NEG POS net36 / NR2HSP_PLL600V3_m18
XI14 net36 NEG POS net73 / IVHSP_PLL600V3_m18
XI8 net4 NEG POS net24 / IVHSP_PLL600V3_m18
XI0 FRIN NEG POS net1 / IVHSP_PLL600V3_m18
XI18 net3 net4 NEG POS / scpllinvsl_PLL600V3_m18
XI19 net1 net3 NEG POS / scpllinvsl_PLL600V3_m18
.ENDS

************************************************************************
* Library Name: SERIAL_LINK_mkm18
* Cell Name:    TIEHI_PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT TIEHI_PLL600V3_m18 NEG POS Y
*.PININFO NEG:I POS:I Y:O
MM0 net09 net09 NEG NEG NHS W=0.3e-6 L=0.18e-6 M=1
MM1 Y net09 POS POS PHS W=1e-6 L=0.18e-6 M=1
.ENDS

************************************************************************
* Library Name: SINT_mkm18
* Cell Name:    FD1HSP_dummy_PLL600V3_m18
* View Name:    cmos_sch
************************************************************************

.SUBCKT FD1HSP_dummy_PLL600V3_m18 CP D NEG POS Q QN
*.PININFO CP:I D:I NEG:I POS:I Q:O QN:O
XI28 NEG POS net106 / TIEHI_PLL600V3_m18
MMN16 Q M4 NEG NEG NHS W=1.42u L=0.18u M=1
MMN11 M4 S1 NEG NEG NHS W=0.80u L=0.18u M=1
MMN103 M1 CN DIN NEG NHS W=0.28u L=0.18u M=1
MMN71 M5N net106 NEG NEG NHS W=0.28u L=0.18u M=1
MMN74 S1 CN M5N NEG NHS W=0.28u L=0.18u M=1
MMN78 M1 CPI M3N NEG NHS W=0.28u L=0.18u M=1
MMN85 M3N M2 NEG NEG NHS W=0.28u L=0.18u M=1
MMN89 M2 M1 NEG NEG NHS W=0.28u L=0.18u M=1
MMN92 S1 CPI MIN NEG NHS W=0.64u L=0.18u M=1
MMN106 DIN D NEG NEG NHS W=0.28u L=0.18u M=1
MMN123 CPI CN NEG NEG NHS W=0.36u L=0.18u M=1
MM0 MIN M1 NEG NEG NHS W=0.64u L=0.18u M=1
MM24 QN S1 NEG NEG NHS W=1.42u L=0.18u M=1
MMN119 CN CP NEG NEG NHS W=0.70u L=0.18u M=1
MMP16 Q M4 POS POS PHS W=2.50u L=0.18u M=1
MMP11 M4 S1 POS POS PHS W=1.10u L=0.18u M=1
MMP127 S1 CN MIP POS PHS W=1.10u L=0.18u M=1
MMP112 M1 CPI DIP POS PHS W=0.56u L=0.18u M=1
MMP72 M5P net106 POS POS PHS W=0.28u L=0.18u M=1
MMP73 S1 CPI M5P POS PHS W=0.28u L=0.18u M=1
MMP76 M1 CN M3P POS PHS W=0.28u L=0.18u M=1
MMP79 M2 M1 POS POS PHS W=0.34u L=0.18u M=1
MMP120 CN CP POS POS PHS W=0.70u L=0.18u M=1
MMP124 CPI CN POS POS PHS W=0.70u L=0.18u M=1
MMP1 MIP M1 POS POS PHS W=1.10u L=0.18u M=1
MM5 QN S1 POS POS PHS W=2.50u L=0.18u M=1
MMP87 M3P M2 POS POS PHS W=0.28u L=0.18u M=1
MMP102 DIP D POS POS PHS W=0.56u L=0.18u M=1
DD16 D POS DP 1.02e-13
DD0 CP POS DP 1.02e-13
.ENDS

************************************************************************
* Library Name: SINT_mkm18
* Cell Name:    scplldivb_PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT scplldivb_PLL600V3_m18 CLK CLKB D DB L NEG POS Q QB T
*.PININFO CLK:I CLKB:I D:I DB:I L:I NEG:I POS:I T:I Q:O QB:O
MM4 QB Q POS POS PHS W=1.62e-6 L=0.18e-6 M=1
MM30 net124 net121 POS POS PHS W=1.62e-6 L=0.18e-6 M=1
MM15 net121 net124 POS POS PHS W=1.62e-6 L=0.18e-6 M=1
MM34 Q QB POS POS PHS W=1.62e-6 L=0.18e-6 M=1
MM13 net135 Q net117 NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM41 net116 DB NEG NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM5 net121 net124 NEG NEG NHS W=0.52e-6 L=0.18e-6 M=1
MM48 Q CLKB net61 NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM43 net110 T NEG NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM19 net111 L net134 NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM14 net135 Q net110 NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM40 net114 DB NEG NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM6 QB Q NEG NEG NHS W=0.52e-6 L=0.18e-6 M=1
MM12 net135 L net116 NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM45 QB CLKB net102 NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM49 Q CLKB net147 NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM51 net61 net121 NEG NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM38 net105 T NEG NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM31 net134 D NEG NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM39 net101 T NEG NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM21 net111 QB net105 NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM28 Q QB NEG NEG NHS W=0.52e-6 L=0.18e-6 M=1
MM32 net108 D NEG NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM20 net111 L net108 NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM22 net111 QB net101 NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM18<0> net124 CLK net135 NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM18<1> net124 CLK net135 NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM11 net135 L net114 NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM37<1> net121 CLK net111 NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM37<0> net121 CLK net111 NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM50 net147 net121 NEG NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM46 net102 net124 NEG NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM27 net124 net121 NEG NEG NHS W=0.52e-6 L=0.18e-6 M=1
MM44 QB CLKB net149 NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM47 net149 net124 NEG NEG NHS W=1.6e-6 L=0.18e-6 M=1
MM42 net117 T NEG NEG NHS W=1.6e-6 L=0.18e-6 M=1
.ENDS

************************************************************************
* Library Name: SERIAL_LINK_mkm18
* Cell Name:    FD4HSP_PLL600V3_m18
* View Name:    cmos_sch
************************************************************************

.SUBCKT FD4HSP_PLL600V3_m18 CP D NEG POS Q QN SD
*.PININFO CP:I D:I NEG:I POS:I SD:I Q:O QN:O
MMN16 Q M4 NEG NEG NHS W=1.42u L=0.18u M=1
MMN11 M4 S1 NEG NEG NHS W=0.80u L=0.18u M=1
MMN103 M1 CN DIN NEG NHS W=0.28u L=0.18u M=1
MMN71 M5N M4 net110 NEG NHS W=0.28u L=0.18u M=1
MMN74 S1 CN M5N NEG NHS W=0.28u L=0.18u M=1
MMN78 M1 CPI M3N NEG NHS W=0.28u L=0.18u M=1
MMN85 M3N M2 NEG NEG NHS W=0.28u L=0.18u M=1
MMN89 M2 M1 net199 NEG NHS W=0.28u L=0.18u M=1
MMN0 MIN M1 MIS NEG NHS W=0.64u L=0.18u M=1
MMN106 DIN D NEG NEG NHS W=0.28u L=0.18u M=1
MMN119 CN CP NEG NEG NHS W=0.70u L=0.18u M=1
MMN123 CPI CN NEG NEG NHS W=0.36u L=0.18u M=1
MMN92 S1 CPI MIN NEG NHS W=0.64u L=0.18u M=1
MMN183 MIS SD NEG NEG NHS W=0.64u L=0.18u M=1
MM7 net110 SD NEG NEG NHS W=0.28u L=0.18u M=1
MM24 QN S1 NEG NEG NHS W=1.42u L=0.18u M=1
MMN83 net199 SD NEG NEG NHS W=0.28u L=0.18u M=1
MMP16 Q M4 POS POS PHS W=2.50u L=0.18u M=1
MMP11 M4 S1 POS POS PHS W=1.10u L=0.18u M=1
MMP190 S1 SD POS POS PHS W=1.10u L=0.18u M=1
MMP112 M1 CPI DIP POS PHS W=0.56u L=0.18u M=1
MMP72 M5P M4 POS POS PHS W=0.28u L=0.18u M=1
MMP73 S1 CPI M5P POS PHS W=0.28u L=0.18u M=1
MMP76 M1 CN M3P POS PHS W=0.28u L=0.18u M=1
MMP79 M2 M1 POS POS PHS W=0.34u L=0.18u M=1
MMP120 CN CP POS POS PHS W=0.70u L=0.18u M=1
MMP124 CPI CN POS POS PHS W=0.70u L=0.18u M=1
MM5 QN S1 POS POS PHS W=2.50u L=0.18u M=1
MMP127 S1 CN MIP POS PHS W=1.10u L=0.18u M=1
MMP1 MIP M1 POS POS PHS W=1.10u L=0.18u M=1
MMP87 M3P M2 POS POS PHS W=0.28u L=0.18u M=1
MMP102 DIP D POS POS PHS W=0.56u L=0.18u M=1
MMP90 M2 SD POS POS PHS W=0.34u L=0.18u M=1
DD16 D POS DP 1.02e-13
DD0 CP POS DP 1.02e-13
DD1 SD POS DP 1.02e-13
.ENDS

************************************************************************
* Library Name: SERIAL_LINK_mkm18
* Cell Name:    IVHSX4_PLL600V3_m18
* View Name:    cmos_sch
************************************************************************

.SUBCKT IVHSX4_PLL600V3_m18 A NEG POS Z
*.PININFO A:I NEG:I POS:I Z:O
MMN1 Z A NEG NEG NHS W=2.84u L=0.18u M=1
MMP1 Z A POS POS PHS W=5.06u L=0.18u M=1
DD7 NEG A DN 1.02e-13
.ENDS

************************************************************************
* Library Name: SERIAL_LINK_mkm18
* Cell Name:    ND4HSP_PLL600V3_m18
* View Name:    cmos_sch
************************************************************************

.SUBCKT ND4HSP_PLL600V3_m18 A B C D NEG POS Z
*.PININFO A:I B:I C:I D:I NEG:I POS:I Z:O
MMN4 net3 D NEG NEG NHS W=1.78u L=0.18u M=1
MMN3 net6 C net3 NEG NHS W=1.78u L=0.18u M=1
MMN2 net9 B net6 NEG NHS W=1.78u L=0.18u M=1
MMN1 Z A net9 NEG NHS W=1.78u L=0.18u M=1
MM22 net22 D NEG NEG NHS W=1.78u L=0.18u M=1
MM21 net25 C net22 NEG NHS W=1.78u L=0.18u M=1
MM20 Z A net31 NEG NHS W=1.78u L=0.18u M=1
MM19 net31 B net25 NEG NHS W=1.78u L=0.18u M=1
MMP1 Z A POS POS PHS W=2.50u L=0.18u M=1
MMP2 Z B POS POS PHS W=2.52u L=0.18u M=1
MMP3 Z C POS POS PHS W=2.52u L=0.18u M=1
MMP4 Z D POS POS PHS W=2.52u L=0.18u M=1
DD38 A POS DP 1.02e-13
DD34 C POS DP 1.02e-13
DD30 B POS DP 1.02e-13
DD24 NEG D DN 1.02e-13
.ENDS

************************************************************************
* Library Name: SERIAL_LINK_mkm18
* Cell Name:    ND3HSP_PLL600V3_m18
* View Name:    cmos_sch
************************************************************************

.SUBCKT ND3HSP_PLL600V3_m18 A B C NEG POS Z
*.PININFO A:I B:I C:I NEG:I POS:I Z:O
MMN3 net3 C NEG NEG NHS W=1.42u L=0.18u M=1
MMN2 net6 B net3 NEG NHS W=1.42u L=0.18u M=1
MMN1 Z A net6 NEG NHS W=1.42u L=0.18u M=1
MM17 net18 C NEG NEG NHS W=1.42u L=0.18u M=1
MM16 net21 B net18 NEG NHS W=1.42u L=0.18u M=1
MM15 Z A net21 NEG NHS W=1.42u L=0.18u M=1
MMP3 Z C POS POS PHS W=2.50u L=0.18u M=1
MMP2 Z B POS POS PHS W=2.52u L=0.18u M=1
MMP1 Z A POS POS PHS W=2.52u L=0.18u M=1
DD24 NEG C DN 1.02e-13
DD25 B POS DP 1.02e-13
DD21 A POS DP 1.02e-13
.ENDS

************************************************************************
* Library Name: SINT_mkm18
* Cell Name:    scplldivid_PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT scplldivid_PLL600V3_m18 CLKINB D0 D1 D2 D3 D4 DIVOUT DIVOUT2 FORCE32 
+ NEG POS RESET SYNCEN
*.PININFO CLKINB:I D0:I D1:I D2:I D3:I D4:I FORCE32:I NEG:I POS:I RESET:I 
*.PININFO SYNCEN:I DIVOUT:O DIVOUT2:O
XI65 net173 net190 NEG POS DIVOUT net233 / FD1HSP_dummy_PLL600V3_m18
XXI58 CLK CLKB net142 net359 LOAD NEG POS Q4 net406 net336 / 
+ scplldivb_PLL600V3_m18
XI57 CLK CLKB net303 net357 LOAD NEG POS Q2 net394 net337 / 
+ scplldivb_PLL600V3_m18
XI58 CLK CLKB net143 net355 LOAD NEG POS Q1 net382 net378 / 
+ scplldivb_PLL600V3_m18
XI56 CLK CLKB net149 net361 LOAD NEG POS Q3 net418 net414 / 
+ scplldivb_PLL600V3_m18
XI59 CLK CLKB net347 net353 LOAD NEG POS Q0 net370 net223 / 
+ scplldivb_PLL600V3_m18
MM5<0> net278 net273 NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM5<1> net278 net273 NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM5<2> net278 net273 NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM5<3> net278 net273 NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM5<4> net278 net273 NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM6<0> CLKB net273 NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM6<1> CLKB net273 NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM6<2> CLKB net273 NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM6<3> CLKB net273 NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM6<4> CLKB net273 NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM7<0> net273 net173 NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM7<1> net273 net173 NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM7<2> net273 net173 NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM7<3> net273 net173 NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM4<0> CLK net278 NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM4<1> CLK net278 NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM4<2> CLK net278 NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM0<0> CLK net278 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM0<1> CLK net278 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM0<2> CLK net278 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM0<3> CLK net278 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM0<4> CLK net278 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM0<5> CLK net278 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM0<6> CLK net278 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM0<7> CLK net278 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM0<8> CLK net278 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM0<9> CLK net278 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM2<0> CLKB net273 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM2<1> CLKB net273 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM2<2> CLKB net273 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM2<3> CLKB net273 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM2<4> CLKB net273 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM2<5> CLKB net273 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM2<6> CLKB net273 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM2<7> CLKB net273 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM2<8> CLKB net273 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM2<9> CLKB net273 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM3<0> net273 net173 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM3<1> net273 net173 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM3<2> net273 net173 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM3<3> net273 net173 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM3<4> net273 net173 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM3<5> net273 net173 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM1<0> net278 net273 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM1<1> net278 net273 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM1<2> net278 net273 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM1<3> net278 net273 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM1<4> net278 net273 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM1<5> net278 net273 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM1<6> net278 net273 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM1<7> net278 net273 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM1<8> net278 net273 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
MM1<9> net278 net273 POS POS PHS W=2.08e-6 L=0.18e-6 M=1
XI50 net173 net138 NEG POS net131 net139 RESB / FD4HSP_PLL600V3_m18
XI49 net173 NEG NEG POS net301 net225 RESB / FD4HSP_PLL600V3_m18
XI39 CLKINB NEG POS net173 / IVHSX4_PLL600V3_m18
XI38 CLKINB NEG POS net173 / IVHSX4_PLL600V3_m18
XI45 net139 NEG POS LOAD / IVHSX4_PLL600V3_m18
XI46 net139 NEG POS LOAD / IVHSX4_PLL600V3_m18
XI33 net274 net146 net175 net123 NEG POS net335 / ND4HSP_PLL600V3_m18
XI32 net274 net146 net175 NEG POS net150 / ND3HSP_PLL600V3_m18
XI18 net136 LOAD NEG POS net378 / NR2HSP_PLL600V3_m18
XI51 net327 net131 NEG POS net197 / NR2HSP_PLL600V3_m18
XI52 net197 net301 NEG POS net190 / NR2HSP_PLL600V3_m18
XI27 net150 LOAD NEG POS net414 / NR2HSP_PLL600V3_m18
XI31 net335 LOAD NEG POS net336 / NR2HSP_PLL600V3_m18
XI48 net245 F32 NEG POS net327 / NR2HSP_PLL600V3_m18
XI16 D1 F32 NEG POS net143 / NR2HSP_PLL600V3_m18
XI29 D4 F32 NEG POS net142 / NR2HSP_PLL600V3_m18
XI22 D2 F32 NEG POS net303 / NR2HSP_PLL600V3_m18
XI25 D3 F32 NEG POS net149 / NR2HSP_PLL600V3_m18
XI44 net335 net95 NEG POS net138 / NR2HSP_PLL600V3_m18
XI21 net271 LOAD NEG POS net337 / NR2HSP_PLL600V3_m18
XI55 net233 net301 NEG POS DIVOUT2 / NR2HSP_PLL600V3_m18
XI36 net139 Q4 NEG POS net2 / ND2HSP_PLL600V3_m18
XI11 D0 net188 NEG POS net347 / ND2HSP_PLL600V3_m18
XI20 net274 net146 NEG POS net271 / ND2HSP_PLL600V3_m18
XI34 net1 NEG POS net95 / IVHSP_PLL600V3_m18
XI17 net143 NEG POS net355 / IVHSP_PLL600V3_m18
XI30 net142 NEG POS net359 / IVHSP_PLL600V3_m18
XI19 net382 NEG POS net146 / IVHSP_PLL600V3_m18
XI10 net188 NEG POS F32 / IVHSP_PLL600V3_m18
XI15 net370 NEG POS net274 / IVHSP_PLL600V3_m18
XI23 net303 NEG POS net357 / IVHSP_PLL600V3_m18
XI14 Q0 NEG POS net136 / IVHSP_PLL600V3_m18
XI24 net394 NEG POS net175 / IVHSP_PLL600V3_m18
XI37 RESET NEG POS RESB / IVHSP_PLL600V3_m18
XI28 net418 NEG POS net123 / IVHSP_PLL600V3_m18
XI35 net2 NEG POS net1 / IVHSP_PLL600V3_m18
XI47 SYNCEN NEG POS net245 / IVHSP_PLL600V3_m18
XI13 LOAD NEG POS net223 / IVHSP_PLL600V3_m18
XI12 net347 NEG POS net353 / IVHSP_PLL600V3_m18
XI9 FORCE32 NEG POS net188 / IVHSP_PLL600V3_m18
XI26 net149 NEG POS net361 / IVHSP_PLL600V3_m18
.ENDS

************************************************************************
* Library Name: SINT_mkm18
* Cell Name:    PLLFILTSUPV2_PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT PLLFILTSUPV2_PLL600V3_m18 FILPOS NEG POS
*.PININFO NEG:I POS:I FILPOS:O
DD1 NEG POS DI 1.00e-12
RR5 FILPOS POS 190.9 $SUB=NEG $[R4] $W=2.1e-6 M=1
RR8 FILPOS POS 190.9 $SUB=NEG $[R4] $W=2.1e-6 M=1
RR11 FILPOS POS 190.9 $SUB=NEG $[R4] $W=2.1e-6 M=1
RR10 FILPOS POS 190.9 $SUB=NEG $[R4] $W=2.1e-6 M=1
RR1 FILPOS POS 190.9 $SUB=NEG $[R4] $W=2.1e-6 M=1
RR7 FILPOS POS 190.9 $SUB=NEG $[R4] $W=2.1e-6 M=1
RR6 FILPOS POS 190.9 $SUB=NEG $[R4] $W=2.1e-6 M=1
RR2 FILPOS POS 190.9 $SUB=NEG $[R4] $W=2.1e-6 M=1
RR3 FILPOS POS 190.9 $SUB=NEG $[R4] $W=2.1e-6 M=1
RR0 FILPOS POS 190.9 $SUB=NEG $[R4] $W=2.1e-6 M=1
RR4 FILPOS POS 190.9 $SUB=NEG $[R4] $W=2.1e-6 M=1
RR9 FILPOS POS 190.9 $SUB=NEG $[R4] $W=2.1e-6 M=1
MM0<1> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<2> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<3> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<4> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<5> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<6> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<7> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<8> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<9> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<10> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<11> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<12> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<13> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<14> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<15> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<16> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<17> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<18> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<19> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<20> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<21> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<22> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<23> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<24> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<25> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<26> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<27> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<28> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<29> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<30> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<31> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<32> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<33> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<34> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<35> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<36> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<37> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<38> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<39> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<40> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<41> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<42> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<43> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<44> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<45> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<46> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<47> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<48> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<49> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<50> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<51> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<52> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<53> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<54> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<55> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<56> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<57> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<58> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<59> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<60> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<61> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<62> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<63> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<64> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<65> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<66> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<67> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<68> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<69> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<70> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<71> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<72> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<73> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<74> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<75> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<76> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<77> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<78> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<79> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<80> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<81> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<82> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<83> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<84> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<85> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<86> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<87> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<88> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<89> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<90> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<91> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<92> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<93> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<94> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<95> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<96> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<97> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<98> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<99> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<100> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<101> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<102> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<103> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<104> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<105> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<106> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<107> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<108> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<109> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<110> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<111> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<112> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<113> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<114> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<115> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<116> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<117> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<118> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<119> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<120> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<121> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<122> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<123> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<124> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<125> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<126> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<127> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<128> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<129> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<130> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<131> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<132> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<133> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<134> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<135> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<136> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<137> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<138> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<139> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<140> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<141> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<142> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<143> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<144> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<145> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<146> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<147> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<148> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<149> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<150> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<151> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<152> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<153> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<154> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<155> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<156> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<157> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<158> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<159> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<160> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<161> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<162> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<163> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<164> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<165> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<166> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<167> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<168> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<169> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<170> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<171> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<172> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<173> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<174> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<175> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<176> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<177> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<178> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<179> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<180> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<181> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<182> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<183> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<184> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<185> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<186> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<187> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<188> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<189> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<190> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<191> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<192> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<193> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<194> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<195> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<196> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<197> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<198> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<199> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<200> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<201> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<202> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<203> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<204> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<205> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<206> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<207> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<208> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<209> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<210> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<211> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<212> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<213> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<214> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<215> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<216> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<217> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<218> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<219> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<220> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<221> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<222> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<223> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<224> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<225> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<226> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<227> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<228> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<229> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<230> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<231> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<232> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<233> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<234> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<235> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<236> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<237> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<238> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<239> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<240> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<241> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<242> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<243> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<244> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<245> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<246> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<247> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<248> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<249> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<250> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<251> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<252> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<253> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<254> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<255> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<256> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<257> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<258> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<259> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<260> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<261> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<262> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<263> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<264> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<265> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<266> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<267> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<268> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<269> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<270> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<271> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<272> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<273> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<274> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<275> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<276> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<277> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<278> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<279> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<280> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<281> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<282> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<283> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<284> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<285> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<286> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<287> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<288> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<289> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<290> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<291> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<292> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<293> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<294> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<295> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<296> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<297> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<298> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<299> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<300> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<301> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<302> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<303> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<304> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<305> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<306> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<307> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<308> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<309> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<310> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<311> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<312> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<313> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<314> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<315> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<316> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<317> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<318> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<319> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<320> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<321> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<322> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<323> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<324> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<325> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<326> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<327> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<328> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<329> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<330> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<331> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<332> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<333> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<334> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<335> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<336> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<337> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<338> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<339> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<340> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<341> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<342> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<343> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<344> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<345> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<346> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<347> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<348> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<349> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<350> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<351> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<352> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<353> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<354> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<355> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<356> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<357> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<358> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<359> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<360> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<361> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<362> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<363> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<364> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<365> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<366> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<367> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<368> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<369> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<370> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<371> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<372> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<373> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<374> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<375> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<376> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<377> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<378> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<379> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<380> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<381> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<382> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<383> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<384> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<385> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<386> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<387> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<388> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<389> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<390> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<391> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<392> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<393> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<394> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<395> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<396> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<397> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<398> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<399> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<400> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<401> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<402> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<403> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<404> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<405> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<406> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<407> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<408> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<409> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<410> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<411> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<412> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<413> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<414> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<415> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<416> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<417> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<418> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<419> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<420> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<421> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<422> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<423> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<424> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<425> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<426> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<427> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<428> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<429> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<430> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<431> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<432> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<433> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<434> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<435> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<436> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<437> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<438> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<439> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<440> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<441> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<442> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<443> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<444> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<445> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<446> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<447> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<448> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<449> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<450> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<451> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<452> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<453> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<454> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<455> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<456> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<457> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<458> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<459> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<460> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<461> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<462> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<463> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<464> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<465> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<466> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<467> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<468> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<469> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<470> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<471> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<472> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<473> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<474> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<475> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<476> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<477> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<478> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<479> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<480> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<481> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<482> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<483> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<484> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<485> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<486> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<487> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<488> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<489> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<490> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<491> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<492> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<493> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<494> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<495> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<496> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<497> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<498> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<499> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<500> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<501> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<502> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<503> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<504> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<505> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<506> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<507> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<508> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<509> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<510> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<511> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<512> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<513> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<514> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<515> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<516> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<517> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<518> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<519> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<520> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<521> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<522> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<523> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<524> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<525> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<526> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<527> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<528> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<529> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<530> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<531> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<532> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<533> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<534> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<535> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<536> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<537> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<538> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<539> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<540> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<541> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<542> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<543> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<544> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<545> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<546> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<547> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<548> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<549> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<550> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<551> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<552> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<553> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<554> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<555> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<556> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<557> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<558> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<559> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<560> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<561> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<562> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<563> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<564> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<565> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<566> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<567> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<568> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<569> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<570> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<571> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<572> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<573> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<574> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<575> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
MM0<576> NEG FILPOS NEG NEG NHS W=9.4e-6 L=4.54e-6 M=1
.ENDS

************************************************************************
* Library Name: SERIAL_LINK_mkm18
* Cell Name:    TIELO_PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT TIELO_PLL600V3_m18 NEG POS Y
*.PININFO NEG:I POS:I Y:O
MM1 net7 net7 POS POS PHS W=0.3e-6 L=0.18e-6 M=1
MM0 Y net7 NEG NEG NHS W=0.56e-6 L=0.18e-6 M=1
.ENDS

************************************************************************
* Library Name: SERIAL_LINK_mkm18
* Cell Name:    MX2HSX2_PLL600V3_m18
* View Name:    cmos_sch
************************************************************************

.SUBCKT MX2HSX2_PLL600V3_m18 A B NEG POS S0 Y
*.PININFO A:I B:I NEG:I POS:I S0:I Y:O
MMP4 net661 net660 net622 POS PHS W=1.10u L=0.18u M=1
MMP3 net661 S0 net18 POS PHS W=1.10u L=0.18u M=1
MMP2 net622 B POS POS PHS W=1.10u L=0.18u M=1
MMP1 net18 A POS POS PHS W=1.10u L=0.18u M=1
MMP22 Y net661 POS POS PHS W=1.24u L=0.18u M=1
MMP28 net660 S0 POS POS PHS W=1.24u L=0.18u M=1
MMN3 net3 B NEG NEG NHS W=0.52u L=0.18u M=1
MMN4 net661 S0 net3 NEG NHS W=0.52u L=0.18u M=1
MMN2 net661 net660 net12 NEG NHS W=0.52u L=0.18u M=1
MMN1 net12 A NEG NEG NHS W=0.52u L=0.18u M=1
MMN23 Y net661 NEG NEG NHS W=0.70u L=0.18u M=1
MMN29 net660 S0 NEG NEG NHS W=0.70u L=0.18u M=1
DD32 S0 POS DP 1.02e-13
DD38 NEG A DN 1.02e-13
DD0 NEG B DN 1.02e-13
.ENDS

************************************************************************
* Library Name: SINT_mkm18
* Cell Name:    pllipmux_PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT pllipmux_PLL600V3_m18 CLKBCKB CLKFDB CLKINB CLKREFB NEG POS TESTCON 
+ TESTI
*.PININFO CLKFDB:I CLKINB:I NEG:I POS:I TESTCON:I TESTI:I CLKBCKB:O CLKREFB:O
XI22 NEG POS TIELO / TIELO_PLL600V3_m18
XI30 TESTI NEG POS net027 / IVHSP_PLL600V3_m18
XI25 CLKINB NEG POS net024 / IVHSP_PLL600V3_m18
XI29 CLKFDB NEG POS net031 / IVHSP_PLL600V3_m18
XI28 net031 net027 NEG POS TESTCON CLKBCKB / MX2HSX2_PLL600V3_m18
XI18 net024 TIELO NEG POS TIELO CLKREFB / MX2HSX2_PLL600V3_m18
.ENDS

************************************************************************
* Library Name: SINT_mkm18
* Cell Name:    scplltfac_PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT scplltfac_PLL600V3_m18 CLKINB DT1 NEG NEWDT1 POS SG1 TM1 TM2
*.PININFO CLKINB:I DT1:I NEG:I POS:I SG1:I TM1:I TM2:I NEWDT1:O
XI36 net174 NEG POS NEWDT1 / IVHSX4_PLL600V3_m18
XI32 TM1 SG1 net93 NEG POS net167 / ND3HSP_PLL600V3_m18
XI17 net163 net144 NEG POS net139 / ND2HSP_PLL600V3_m18
XI16 net73 net149 NEG POS net144 / ND2HSP_PLL600V3_m18
XI34 net230 net167 NEG POS net169 / ND2HSP_PLL600V3_m18
XI35 net169 net173 NEG POS net174 / ND2HSP_PLL600V3_m18
XI18 net114 net139 NEG POS net163 / ND2HSP_PLL600V3_m18
XI33 net89 net163 NEG POS net173 / ND2HSP_PLL600V3_m18
XI15 net105 net177 NEG POS net114 / ND2HSP_PLL600V3_m18
XI20 net210 NEG POS net73 / IVHSP_PLL600V3_m18
XI4 net20 NEG POS net177 / IVHSP_PLL600V3_m18
XI1 net167 NEG POS net89 / IVHSP_PLL600V3_m18
XI25 net19 NEG POS net16 / IVHSP_PLL600V3_m18
XI3 net230 NEG POS net105 / IVHSP_PLL600V3_m18
XI2 DT1 NEG POS net230 / IVHSP_PLL600V3_m18
XI13 net9 NEG POS net20 / IVHSP_PLL600V3_m18
XI5 net105 NEG POS net8 / IVHSP_PLL600V3_m18
XI26 net10 NEG POS net19 / IVHSP_PLL600V3_m18
XI23 net18 NEG POS net17 / IVHSP_PLL600V3_m18
XI22 net15 NEG POS net18 / IVHSP_PLL600V3_m18
XI19 CLKINB NEG POS net210 / IVHSP_PLL600V3_m18
XI21 net17 NEG POS net149 / IVHSP_PLL600V3_m18
XI24 net16 NEG POS net15 / IVHSP_PLL600V3_m18
XI30 net13 NEG POS net14 / IVHSP_PLL600V3_m18
XI29 net14 NEG POS net12 / IVHSP_PLL600V3_m18
XI31 net73 NEG POS net13 / IVHSP_PLL600V3_m18
XI28 net12 NEG POS net11 / IVHSP_PLL600V3_m18
XI27 net11 NEG POS net10 / IVHSP_PLL600V3_m18
XI14 net7 NEG POS net9 / IVHSP_PLL600V3_m18
XI6 net8 NEG POS net2 / IVHSP_PLL600V3_m18
XI12 net6 NEG POS net7 / IVHSP_PLL600V3_m18
XI11 net5 NEG POS net6 / IVHSP_PLL600V3_m18
XI10 net4 NEG POS net5 / IVHSP_PLL600V3_m18
XI9 net3 NEG POS net4 / IVHSP_PLL600V3_m18
XI8 net1 NEG POS net3 / IVHSP_PLL600V3_m18
XI7 net2 NEG POS net1 / IVHSP_PLL600V3_m18
XI0 TM2 NEG POS net93 / IVHSP_PLL600V3_m18
.ENDS

************************************************************************
* Library Name: SERIAL_LINK_mkm18
* Cell Name:    AN3HSP_PLL600V3_m18
* View Name:    cmos_sch
************************************************************************

.SUBCKT AN3HSP_PLL600V3_m18 A B C NEG POS Z
*.PININFO A:I B:I C:I NEG:I POS:I Z:O
MMP4 Z net4 POS POS PHS W=2.50u L=0.18u M=1
MMP3 net4 C POS POS PHS W=0.62u L=0.18u M=1
MMP2 net4 B POS POS PHS W=0.62u L=0.18u M=1
MMP1 net4 A POS POS PHS W=0.62u L=0.18u M=1
MMN4 Z net4 NEG NEG NHS W=1.42u L=0.18u M=1
MMN3 net6 C NEG NEG NHS W=0.62u L=0.18u M=1
MMN2 net9 B net6 NEG NHS W=0.62u L=0.18u M=1
MMN1 net4 A net9 NEG NHS W=0.62u L=0.18u M=1
DD5 NEG B DN 1.02e-13
DD29 C POS DP 1.02e-13
DD21 A POS DP 1.02e-13
.ENDS

************************************************************************
* Library Name: SERIAL_LINK_mkm18
* Cell Name:    OR3HSP_PLL600V3_m18
* View Name:    cmos_sch
************************************************************************

.SUBCKT OR3HSP_PLL600V3_m18 A B C NEG POS Z
*.PININFO A:I B:I C:I NEG:I POS:I Z:O
MMP5 Z net19 POS POS PHS W=2.50u L=0.18u M=1
MMP4 net19 A net6 POS PHS W=1.54u L=0.18u M=1
MMP3 net6 B net9 POS PHS W=1.54u L=0.18u M=1
MMP2 net9 C POS POS PHS W=1.54u L=0.18u M=1
MMN5 Z net19 NEG NEG NHS W=1.44u L=0.18u M=1
MMN2 net19 C NEG NEG NHS W=0.34u L=0.18u M=1
MMN3 net19 B NEG NEG NHS W=0.34u L=0.18u M=1
MMN4 net19 A NEG NEG NHS W=0.34u L=0.18u M=1
DD29 B POS DP 1.02e-13
DD1 NEG A DN 1.02e-13
DD23 NEG C DN 1.02e-13
.ENDS

************************************************************************
* Library Name: SERIAL_LINK_mkm18
* Cell Name:    F_EOHSP_PLL600V3_m18
* View Name:    cmos_sch
************************************************************************

.SUBCKT F_EOHSP_PLL600V3_m18 A B NEG POS Z
*.PININFO A:I B:I NEG:I POS:I Z:O
MM22 net84 net80 net59 POS PHS W=1.66u L=0.18u M=1
MM23 net59 net68 POS POS PHS W=1.66u L=0.18u M=1
MM15 net84 B net80 POS PHS W=0.28u L=0.18u M=1
MM16 net84 A net68 POS PHS W=0.28u L=0.18u M=1
MM7 Z net84 POS POS PHS W=2.82u L=0.18u M=1
MM6 net68 B POS POS PHS W=1.70u L=0.18u M=1
MM5 net80 A POS POS PHS W=1.72u L=0.18u M=1
MM17 net84 net80 net68 NEG NHS W=0.66u L=0.18u M=1
MM10 Z net84 NEG NEG NHS W=1.94u L=0.18u M=1
MM9 net68 B NEG NEG NHS W=1.58u L=0.18u M=1
MM14 net84 net68 net80 NEG NHS W=0.66u L=0.18u M=1
MM8 net80 A NEG NEG NHS W=1.60u L=0.18u M=1
DD0 A POS DP 1.02e-13
DD1 NEG B DN 1.02e-13
.ENDS

************************************************************************
* Library Name: SERIAL_LINK_mkm18
* Cell Name:    NR3HSP_PLL600V3_m18
* View Name:    cmos_sch
************************************************************************

.SUBCKT NR3HSP_PLL600V3_m18 A B C NEG POS Z
*.PININFO A:I B:I C:I NEG:I POS:I Z:O
MMP1 net14 net13 POS POS PHS W=1.24u L=0.18u M=1
MM12 Z net14 POS POS PHS W=2.50u L=0.18u M=1
MMP3 net13 A net33 POS PHS W=1.54u L=0.18u M=1
MM13 net39 C POS POS PHS W=1.54u L=0.18u M=1
MMP2 net33 B net39 POS PHS W=1.54u L=0.18u M=1
MM14 net13 C NEG NEG NHS W=0.34u L=0.18u M=1
MMN1 net14 net13 NEG NEG NHS W=0.70u L=0.18u M=1
MM11 Z net14 NEG NEG NHS W=1.42u L=0.18u M=1
MMN3 net13 A NEG NEG NHS W=0.34u L=0.18u M=1
MMN2 net13 B NEG NEG NHS W=0.34u L=0.18u M=1
DD33 B POS DP 1.02e-13
DD20 C POS DP 1.02e-13
DD29 NEG A DN 1.02e-13
.ENDS

************************************************************************
* Library Name: SERIAL_LINK_mkm18
* Cell Name:    OR2HSP_PLL600V3_m18
* View Name:    cmos_sch
************************************************************************

.SUBCKT OR2HSP_PLL600V3_m18 A B NEG POS Z
*.PININFO A:I B:I NEG:I POS:I Z:O
MMN3 Z net13 NEG NEG NHS W=1.44u L=0.18u M=1
MMN2 net13 A NEG NEG NHS W=0.34u L=0.18u M=1
MMN1 net13 B NEG NEG NHS W=0.34u L=0.18u M=1
MMP3 Z net13 POS POS PHS W=2.50u L=0.18u M=1
MMP2 net13 A net6 POS PHS W=1.10u L=0.18u M=1
MMP1 net6 B POS POS PHS W=1.10u L=0.18u M=1
DD17 B POS DP 1.02e-13
DD19 NEG A DN 1.02e-13
.ENDS

************************************************************************
* Library Name: SERIAL_LINK_mkm18
* Cell Name:    AN2HSP_PLL600V3_m18
* View Name:    cmos_sch
************************************************************************

.SUBCKT AN2HSP_PLL600V3_m18 A B NEG POS Z
*.PININFO A:I B:I NEG:I POS:I Z:O
MMP2 net4 B POS POS PHS W=0.62u L=0.18u M=1
MMP3 Z net4 POS POS PHS W=2.50u L=0.18u M=1
MMP1 net4 A POS POS PHS W=0.62u L=0.18u M=1
MMN3 Z net4 NEG NEG NHS W=1.42u L=0.18u M=1
MMN2 net6 B NEG NEG NHS W=0.52u L=0.18u M=1
MMN1 net4 A net6 NEG NHS W=0.52u L=0.18u M=1
DD26 B POS DP 1.02e-13
DD20 NEG A DN 1.02e-13
.ENDS

************************************************************************
* Library Name: SINT_mkm18
* Cell Name:    scplltogd_PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT scplltogd_PLL600V3_m18 IN NEG OUT POS
*.PININFO IN:I NEG:I POS:I OUT:O
XI12 net8 net13 NEG POS OUT / F_EOHSP_PLL600V3_m18
XI1 net8 NEG POS net10 / IVHSP_PLL600V3_m18
XI9 net2 NEG POS net1 / IVHSP_PLL600V3_m18
XI6 net7 NEG POS net4 / IVHSP_PLL600V3_m18
XI2 net10 NEG POS net9 / IVHSP_PLL600V3_m18
XI3 net9 NEG POS net6 / IVHSP_PLL600V3_m18
XI5 net5 NEG POS net7 / IVHSP_PLL600V3_m18
XI4 net6 NEG POS net5 / IVHSP_PLL600V3_m18
XI0 IN NEG POS net8 / IVHSP_PLL600V3_m18
XI7 net4 NEG POS net3 / IVHSP_PLL600V3_m18
XI8 net3 NEG POS net2 / IVHSP_PLL600V3_m18
XI10 net1 NEG POS net13 / IVHSP_PLL600V3_m18
.ENDS

************************************************************************
* Library Name: SINT_mkm18
* Cell Name:    scplltcon_PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT scplltcon_PLL600V3_m18 CHPTEST CLKFDB DIVRES DT1 ENB FORCE32 NEG PD 
+ PDANA POS SG1 TM1 TM2 VCOTEST
*.PININFO CLKFDB:I ENB:I NEG:I PD:I POS:I SG1:I TM1:I TM2:I CHPTEST:O DIVRES:O 
*.PININFO DT1:O FORCE32:O PDANA:O VCOTEST:O
XI35 TM1 TM2B SG1B NEG POS VCOTEST / AN3HSP_PLL600V3_m18
XI34 TOGTM1 TOGTM2 TOGSG1 NEG POS CRES / OR3HSP_PLL600V3_m18
XI36 CRES net65 PDANA NEG POS DIVRES / OR3HSP_PLL600V3_m18
XI33 TM2B SG1 NEG POS net16 / F_EOHSP_PLL600V3_m18
XI32 TM1 TM2 PDB NEG POS MODE1PD / NR3HSP_PLL600V3_m18
XI30 net71 net146 VCOTEST NEG POS net72 / ND3HSP_PLL600V3_m18
XI28 net149 NEG POS DT1 / IVHSX4_PLL600V3_m18
XI17 MODE2 MODE1PD NEG POS PDANA / OR2HSP_PLL600V3_m18
XI31 net72 net69 NEG POS net71 / ND2HSP_PLL600V3_m18
XI14 CLKFDB TM1 NEG POS net69 / ND2HSP_PLL600V3_m18
XI10 TM1 TM2 NEG POS CHPTEST / AN2HSP_PLL600V3_m18
XI11 TM1 SG1 NEG POS net44 / AN2HSP_PLL600V3_m18
XI13 TM1B TM2 NEG POS MODE2 / AN2HSP_PLL600V3_m18
XI9 TM1 net16 NEG POS FORCE32 / AN2HSP_PLL600V3_m18
XI8 net44 NEG TOGSG1 POS / scplltogd_PLL600V3_m18
XI7 TM2 NEG TOGTM2 POS / scplltogd_PLL600V3_m18
XXI19 TM1 NEG TOGTM1 POS / scplltogd_PLL600V3_m18
XI15 PD ENB NEG POS PDB / NR2HSP_PLL600V3_m18
XI26 DIVRES NEG POS net146 / IVHSP_PLL600V3_m18
XI25 net10 NEG POS net65 / IVHSP_PLL600V3_m18
XI19 net67 NEG POS net11 / IVHSP_PLL600V3_m18
XI12 TM1 NEG POS TM1B / IVHSP_PLL600V3_m18
XI5 TM2 NEG POS TM2B / IVHSP_PLL600V3_m18
XI24 net3 NEG POS net10 / IVHSP_PLL600V3_m18
XI20 net11 NEG POS net2 / IVHSP_PLL600V3_m18
XI27 net71 NEG POS net149 / IVHSP_PLL600V3_m18
XI23 net1 NEG POS net4 / IVHSP_PLL600V3_m18
XI22 net4 NEG POS net3 / IVHSP_PLL600V3_m18
XI21 net2 NEG POS net1 / IVHSP_PLL600V3_m18
XI18 CRES NEG POS net67 / IVHSP_PLL600V3_m18
XI4 SG1 NEG POS SG1B / IVHSP_PLL600V3_m18
.ENDS

************************************************************************
* Library Name: SINT_mkm18
* Cell Name:    scpllphdet_PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT scpllphdet_PLL600V3_m18 CLKBCKB CLKREFB DN DNB MONBCK MONREF NEG 
+ PHDDNB PHDUPB POS UP UPB
*.PININFO CLKBCKB:I CLKREFB:I NEG:I POS:I DN:O DNB:O MONBCK:O MONREF:O 
*.PININFO PHDDNB:O PHDUPB:O UP:O UPB:O
XI59 net41 NEG POS CUP / IVHSX4_PLL600V3_m18
XI58 net1 NEG POS CDN / IVHSX4_PLL600V3_m18
XI55 net32 net22 net70 NEG POS net41 / ND3HSP_PLL600V3_m18
XI56 net56 net46 net32 NEG POS net1 / ND3HSP_PLL600V3_m18
XI39 CLKREFB NEG POS MONREF / IVHSP_PLL600V3_m18
XI42 net43 NEG POS DN / IVHSP_PLL600V3_m18
XI47 CUP NEG POS net35 / IVHSP_PLL600V3_m18
XI46 CUP NEG POS net42 / IVHSP_PLL600V3_m18
XI51 net3 NEG POS UPB / IVHSP_PLL600V3_m18
XI49 net42 NEG POS net3 / IVHSP_PLL600V3_m18
XI43 net36 NEG POS net2 / IVHSP_PLL600V3_m18
XI50 CUP NEG POS PHDUPB / IVHSP_PLL600V3_m18
XI48 net35 NEG POS UP / IVHSP_PLL600V3_m18
XI52 net2 NEG POS DNB / IVHSP_PLL600V3_m18
XI54 CLKBCKB NEG POS MONBCK / IVHSP_PLL600V3_m18
XI45 CDN NEG POS net43 / IVHSP_PLL600V3_m18
XI44 CDN NEG POS net36 / IVHSP_PLL600V3_m18
XI41 CDN NEG POS PHDDNB / IVHSP_PLL600V3_m18
XI37 net66 net70 NEG POS net22 / ND2HSP_PLL600V3_m18
XI36 net32 net22 NEG POS net66 / ND2HSP_PLL600V3_m18
XI35 CDN CUP NEG POS net32 / ND2HSP_PLL600V3_m18
XI38 net41 CLKBCKB NEG POS net70 / ND2HSP_PLL600V3_m18
XI34 CLKREFB net1 NEG POS net56 / ND2HSP_PLL600V3_m18
XI33 net46 net32 NEG POS net44 / ND2HSP_PLL600V3_m18
XI32 net56 net44 NEG POS net46 / ND2HSP_PLL600V3_m18
.ENDS

************************************************************************
* Library Name: SERIAL_LINK_mkm18
* Cell Name:    NR2HS_PLL600V3_m18
* View Name:    cmos_sch
************************************************************************

.SUBCKT NR2HS_PLL600V3_m18 A B NEG POS Z
*.PININFO A:I B:I NEG:I POS:I Z:O
MMP2 Z A net3 POS PHS W=2.30u L=0.18u M=1
MMP1 net3 B POS POS PHS W=2.30u L=0.18u M=1
MMN1 Z B NEG NEG NHS W=0.88u L=0.18u M=1
MMN2 Z A NEG NEG NHS W=0.88u L=0.18u M=1
DD15 NEG A DN 1.02e-13
DD0 NEG B DN 1.02e-13
.ENDS

************************************************************************
* Library Name: SINT_mkm18
* Cell Name:    scplllkdet_PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT scplllkdet_PLL600V3_m18 LKDET MONBCK MONREF NEG PD PHDDNB PHDUPB POS
*.PININFO MONBCK:I MONREF:I NEG:I PD:I PHDDNB:I PHDUPB:I POS:I LKDET:O
DD1 NEG POS DI 1.00e-12
XI101 PD NEG POS S / IVHSX4_PLL600V3_m18
XI112 net098 NEG POS net093 / IVHSP_PLL600V3_m18
XI114 net093 NEG POS net094 / IVHSP_PLL600V3_m18
XI113 net097 NEG POS net098 / IVHSP_PLL600V3_m18
XI111 net0110 NEG POS net0106 / IVHSP_PLL600V3_m18
XI109 net0106 NEG POS net097 / IVHSP_PLL600V3_m18
XI103 net065 NEG POS net0141 / IVHSP_PLL600V3_m18
XI108 net0117 NEG POS net0133 / IVHSP_PLL600V3_m18
XI115 net094 NEG POS net042 / IVHSP_PLL600V3_m18
XI110 PHDDNB NEG POS net0110 / IVHSP_PLL600V3_m18
XI107 PHDUPB NEG POS net0125 / IVHSP_PLL600V3_m18
XI106 net0125 NEG POS net0117 / IVHSP_PLL600V3_m18
XI96 net074 NEG POS LKDET / IVHSP_PLL600V3_m18
XI95 net091 NEG POS net074 / IVHSP_PLL600V3_m18
XI105 net066 NEG POS net065 / IVHSP_PLL600V3_m18
XI104 net0133 NEG POS net066 / IVHSP_PLL600V3_m18
XI102 net0141 NEG POS net046 / IVHSP_PLL600V3_m18
XI91 A B NEG POS XR / NR2HS_PLL600V3_m18
XI92 net079 net0134 NEG POS net0137 net0134 XR / FD4HSP_PLL600V3_m18
XI98 MONREF net046 NEG POS A net105 S / FD4HSP_PLL600V3_m18
XI100 net0137 net0127 NEG POS net0130 net0127 XR / FD4HSP_PLL600V3_m18
XI99 net086 net076 NEG POS net079 net076 XR / FD4HSP_PLL600V3_m18
XI84 net051 net041 NEG POS net044 net041 XR / FD4HSP_PLL600V3_m18
XI97 MONBCK net042 NEG POS B net98 S / FD4HSP_PLL600V3_m18
XI86 net037 net027 NEG POS net030 net027 XR / FD4HSP_PLL600V3_m18
XI85 net044 net034 NEG POS net037 net034 XR / FD4HSP_PLL600V3_m18
XI89 net079 NEG NEG POS net054 net091 XR / FD4HSP_PLL600V3_m18
XI87 net030 net083 NEG POS net086 net083 XR / FD4HSP_PLL600V3_m18
XI83 MONBCK net048 NEG POS net051 net048 XR / FD4HSP_PLL600V3_m18
.ENDS

************************************************************************
* Library Name: SINT_mkm18
* Cell Name:    scpllchgpmp_PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT scpllchgpmp_PLL600V3_m18 BUFOUT CHP0 CHP1 CHP2 CHP3 CHP4 CHPOUT DN DNB 
+ IREF NEG PDANA POS UP UPB VCOTEST
*.PININFO CHP0:I CHP1:I CHP2:I CHP3:I CHP4:I DN:I DNB:I NEG:I PDANA:I POS:I 
*.PININFO UP:I UPB:I VCOTEST:I CHPOUT:O IREF:O BUFOUT:B
DD1 NEG POS DI 1.00e-12
RR9 net13 net11 814 $SUB=POS $[R4] $W=2.1e-6 M=1
RR1 POS net6 814 $SUB=POS $[R4] $W=2.1e-6 M=1
RR8 net12 net13 814 $SUB=POS $[R4] $W=2.1e-6 M=1
RR7 net8 net12 814 $SUB=POS $[R4] $W=2.1e-6 M=1
RR12 net_258 net10 814 $SUB=POS $[R4] $W=2.1e-6 M=1
RR5 net7 net3 814 $SUB=POS $[R4] $W=2.1e-6 M=1
RR10 net9 net11 814 $SUB=POS $[R4] $W=2.1e-6 M=1
RR3 net5 net2 814 $SUB=POS $[R4] $W=2.1e-6 M=1
RR11 net10 net9 814 $SUB=POS $[R4] $W=2.1e-6 M=1
RR6 net8 net7 814 $SUB=POS $[R4] $W=2.1e-6 M=1
RR2 net6 net5 814 $SUB=POS $[R4] $W=2.1e-6 M=1
RR4 net3 net2 814 $SUB=POS $[R4] $W=2.1e-6 M=1
MM74<0> net79 CHPOUT net46 POS PHS W=10e-6 L=500e-9 M=1
MM74<1> net79 CHPOUT net46 POS PHS W=10e-6 L=500e-9 M=1
MM74<2> net79 CHPOUT net46 POS PHS W=10e-6 L=500e-9 M=1
MM74<3> net79 CHPOUT net46 POS PHS W=10e-6 L=500e-9 M=1
MM74<4> net79 CHPOUT net46 POS PHS W=10e-6 L=500e-9 M=1
MM74<5> net79 CHPOUT net46 POS PHS W=10e-6 L=500e-9 M=1
MM74<6> net79 CHPOUT net46 POS PHS W=10e-6 L=500e-9 M=1
MM74<7> net79 CHPOUT net46 POS PHS W=10e-6 L=500e-9 M=1
MM45 CHP0INT CHP0 POS POS PHS W=4e-6 L=1e-6 M=1
MM48<3> net_191 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM48<2> net_191 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM48<1> net_191 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM48<0> net_191 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM37 net_282 PD POS POS PHS W=1e-6 L=8e-6 M=1
MM67 CHPOUT UPB net_236 POS PHS W=1e-6 L=180e-9 M=1
MM56 net_310 CHP0INT net_167 POS PHS W=1e-6 L=340e-9 M=1
MM36 PDB PD POS POS PHS W=4e-6 L=1e-6 M=1
MM40<1> net_262 net_258 POS POS PHS W=4e-6 L=1e-6 M=1
MM40<0> net_262 net_258 POS POS PHS W=4e-6 L=1e-6 M=1
MM53 CHP3INT CHP3 POS POS PHS W=4e-6 L=1e-6 M=1
MM55 CHP1INT CHP1 POS POS PHS W=4e-6 L=1e-6 M=1
MM54 CHP2INT CHP2 POS POS PHS W=4e-6 L=1e-6 M=1
MM63 net_273 PDB POS POS PHS W=4e-6 L=1e-6 M=1
MM47<1> net_188 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM47<0> net_188 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM57 net_310 CHP1INT net_188 POS PHS W=1e-6 L=340e-9 M=1
MM66 net_236 net_297 net_170 POS PHS W=6e-6 L=500e-9 M=1
MM50<15> net_197 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM50<14> net_197 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM50<13> net_197 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM50<12> net_197 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM50<11> net_197 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM50<10> net_197 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM50<9> net_197 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM50<8> net_197 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM50<7> net_197 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM50<6> net_197 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM50<5> net_197 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM50<4> net_197 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM50<3> net_197 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM50<2> net_197 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM50<1> net_197 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM50<0> net_197 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM51<9> net1 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM51<8> net1 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM51<7> net1 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM51<6> net1 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM51<5> net1 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM51<4> net1 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM51<3> net1 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM51<2> net1 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM51<1> net1 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM51<0> net1 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM62<3> net_173 net_273 POS POS PHS W=10e-6 L=3e-6 M=1
MM62<2> net_173 net_273 POS POS PHS W=10e-6 L=3e-6 M=1
MM62<1> net_173 net_273 POS POS PHS W=10e-6 L=3e-6 M=1
MM62<0> net_173 net_273 POS POS PHS W=10e-6 L=3e-6 M=1
MM59 net_310 CHP3INT net_194 POS PHS W=1e-6 L=340e-9 M=1
MM58 net_310 CHP2INT net_191 POS PHS W=1e-6 L=340e-9 M=1
MM61<3> net_170 net_273 POS POS PHS W=10e-6 L=3e-6 M=1
MM61<2> net_170 net_273 POS POS PHS W=10e-6 L=3e-6 M=1
MM61<1> net_170 net_273 POS POS PHS W=10e-6 L=3e-6 M=1
MM61<0> net_170 net_273 POS POS PHS W=10e-6 L=3e-6 M=1
MM60 net_310 CHP4INT net_197 POS PHS W=1e-6 L=340e-9 M=1
MM69<0> net38 net38 POS POS PHS W=4e-6 L=2e-6 M=1
MM69<1> net38 net38 POS POS PHS W=4e-6 L=2e-6 M=1
MM69<2> net38 net38 POS POS PHS W=4e-6 L=2e-6 M=1
MM69<3> net38 net38 POS POS PHS W=4e-6 L=2e-6 M=1
MM42 net512 net294 POS POS PHS W=4e-6 L=1e-6 M=1
MM52 CHP4INT CHP4 POS POS PHS W=4e-6 L=1e-6 M=1
MM65 net_273 net_297 net_173 POS PHS W=6e-6 L=500e-9 M=1
MM41<3> net294 net294 POS POS PHS W=4e-6 L=1e-6 M=1
MM41<2> net294 net294 POS POS PHS W=4e-6 L=1e-6 M=1
MM41<1> net294 net294 POS POS PHS W=4e-6 L=1e-6 M=1
MM41<0> net294 net294 POS POS PHS W=4e-6 L=1e-6 M=1
MM35 PD net4 POS POS PHS W=4e-6 L=1e-6 M=1
MM44 IREF net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM46 net_167 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM49<7> net_194 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM49<6> net_194 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM49<5> net_194 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM49<4> net_194 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM49<3> net_194 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM49<2> net_194 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM49<1> net_194 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM49<0> net_194 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM70<0> BUFOUT net38 POS POS PHS W=4e-6 L=2e-6 M=1
MM70<1> BUFOUT net38 POS POS PHS W=4e-6 L=2e-6 M=1
MM70<2> BUFOUT net38 POS POS PHS W=4e-6 L=2e-6 M=1
MM70<3> BUFOUT net38 POS POS PHS W=4e-6 L=2e-6 M=1
MM70<4> BUFOUT net38 POS POS PHS W=4e-6 L=2e-6 M=1
MM70<5> BUFOUT net38 POS POS PHS W=4e-6 L=2e-6 M=1
MM70<6> BUFOUT net38 POS POS PHS W=4e-6 L=2e-6 M=1
MM70<7> BUFOUT net38 POS POS PHS W=4e-6 L=2e-6 M=1
MM70<8> BUFOUT net38 POS POS PHS W=4e-6 L=2e-6 M=1
MM70<9> BUFOUT net38 POS POS PHS W=4e-6 L=2e-6 M=1
MM70<10> BUFOUT net38 POS POS PHS W=4e-6 L=2e-6 M=1
MM70<11> BUFOUT net38 POS POS PHS W=4e-6 L=2e-6 M=1
MM70<12> BUFOUT net38 POS POS PHS W=4e-6 L=2e-6 M=1
MM70<13> BUFOUT net38 POS POS PHS W=4e-6 L=2e-6 M=1
MM70<14> BUFOUT net38 POS POS PHS W=4e-6 L=2e-6 M=1
MM70<15> BUFOUT net38 POS POS PHS W=4e-6 L=2e-6 M=1
MM75<0> net32 BUFOUT net46 POS PHS W=10e-6 L=500e-9 M=1
MM75<1> net32 BUFOUT net46 POS PHS W=10e-6 L=500e-9 M=1
MM75<2> net32 BUFOUT net46 POS PHS W=10e-6 L=500e-9 M=1
MM75<3> net32 BUFOUT net46 POS PHS W=10e-6 L=500e-9 M=1
MM75<4> net32 BUFOUT net46 POS PHS W=10e-6 L=500e-9 M=1
MM75<5> net32 BUFOUT net46 POS PHS W=10e-6 L=500e-9 M=1
MM75<6> net32 BUFOUT net46 POS PHS W=10e-6 L=500e-9 M=1
MM75<7> net32 BUFOUT net46 POS PHS W=10e-6 L=500e-9 M=1
MM71<0> IBIAS IBIAS POS POS PHS W=5e-6 L=1e-6 M=1
MM71<1> IBIAS IBIAS POS POS PHS W=5e-6 L=1e-6 M=1
MM71<2> IBIAS IBIAS POS POS PHS W=5e-6 L=1e-6 M=1
MM71<3> IBIAS IBIAS POS POS PHS W=5e-6 L=1e-6 M=1
MM34 net_233 VCOTEST POS POS PHS W=4e-6 L=1e-6 M=1
MM72<0> net46 IBIAS POS POS PHS W=5e-6 L=1e-6 M=1
MM72<1> net46 IBIAS POS POS PHS W=5e-6 L=1e-6 M=1
MM72<2> net46 IBIAS POS POS PHS W=5e-6 L=1e-6 M=1
MM72<3> net46 IBIAS POS POS PHS W=5e-6 L=1e-6 M=1
MM72<4> net46 IBIAS POS POS PHS W=5e-6 L=1e-6 M=1
MM72<5> net46 IBIAS POS POS PHS W=5e-6 L=1e-6 M=1
MM38 net4 PDANA net_233 POS PHS W=4e-6 L=1e-6 M=1
MM43<9> net_261 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM43<8> net_261 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM43<7> net_261 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM43<6> net_261 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM43<5> net_261 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM43<4> net_261 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM43<3> net_261 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM43<2> net_261 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM43<1> net_261 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM43<0> net_261 net_261 POS POS PHS W=1e-6 L=4.84e-6 M=1
MM68 BUFOUT UP net_236 POS PHS W=1e-6 L=180e-9 M=1
MM64 net_297 net_297 POS POS PHS W=3e-6 L=7e-6 M=1
MM14 CHP1INT CHP1 NEG NEG NHS W=4e-6 L=1e-6 M=1
MM15 CHP2INT CHP2 NEG NEG NHS W=4e-6 L=1e-6 M=1
MM17 CHP4INT CHP4 NEG NEG NHS W=4e-6 L=1e-6 M=1
MM16 CHP3INT CHP3 NEG NEG NHS W=4e-6 L=1e-6 M=1
MM12 IBIAS net512 NEG NEG NHS W=4e-6 L=2e-6 M=1
MM29 BUFOUT DNB net_267 NEG NHS W=1e-6 L=180e-9 M=1
MM26<1> net_327 net_310 NEG NEG NHS W=7.5e-6 L=3e-6 M=1
MM26<0> net_327 net_310 NEG NEG NHS W=7.5e-6 L=3e-6 M=1
MM23<1> net_285 net_310 NEG NEG NHS W=7.5e-6 L=3e-6 M=1
MM23<0> net_285 net_310 NEG NEG NHS W=7.5e-6 L=3e-6 M=1
MM10 net512 PD NEG NEG NHS W=4e-6 L=1e-6 M=1
MM20 net_310 net1 net_312 NEG NHS W=3e-6 L=500e-9 M=1
MM8<3> net_262 net_262 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM8<2> net_262 net_262 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM8<1> net_262 net_262 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM8<0> net_262 net_262 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM25 net_310 PD NEG NEG NHS W=4e-6 L=1e-6 M=1
MM6<7> net_258 net512 NEG NEG NHS W=4e-6 L=2e-6 M=1
MM6<6> net_258 net512 NEG NEG NHS W=4e-6 L=2e-6 M=1
MM6<5> net_258 net512 NEG NEG NHS W=4e-6 L=2e-6 M=1
MM6<4> net_258 net512 NEG NEG NHS W=4e-6 L=2e-6 M=1
MM6<3> net_258 net512 NEG NEG NHS W=4e-6 L=2e-6 M=1
MM6<2> net_258 net512 NEG NEG NHS W=4e-6 L=2e-6 M=1
MM6<1> net_258 net512 NEG NEG NHS W=4e-6 L=2e-6 M=1
MM6<0> net_258 net512 NEG NEG NHS W=4e-6 L=2e-6 M=1
MM7 net512 net_262 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM21<1> net_312 net_310 NEG NEG NHS W=7.5e-6 L=3e-6 M=1
MM21<0> net_312 net_310 NEG NEG NHS W=7.5e-6 L=3e-6 M=1
MM24 net_273 net1 net_285 NEG NHS W=3e-6 L=500e-9 M=1
MM27 net_267 net1 net_327 NEG NHS W=3e-6 L=500e-9 M=1
MM11 net_261 net512 NEG NEG NHS W=4e-6 L=2e-6 M=1
MM9 net294 net512 NEG NEG NHS W=4e-6 L=2e-6 M=1
MM13 CHP0INT CHP0 NEG NEG NHS W=4e-6 L=1e-6 M=1
MM19 net1 net1 NEG NEG NHS W=2e-6 L=7.94e-6 M=1
MM22 net_297 net_310 NEG NEG NHS W=4e-6 L=5.94e-6 M=1
MM39<1> POS net_282 net512 NEG NHS W=1e-6 L=4e-6 M=1
MM39<0> POS net_282 net512 NEG NHS W=1e-6 L=4e-6 M=1
MM28 CHPOUT DN net_267 NEG NHS W=1e-6 L=180e-9 M=1
MM30<0> BUFOUT net79 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM30<1> BUFOUT net79 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM30<2> BUFOUT net79 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM30<3> BUFOUT net79 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM30<4> BUFOUT net79 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM30<5> BUFOUT net79 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM30<6> BUFOUT net79 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM30<7> BUFOUT net79 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM32 net32 net32 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM33<0> net38 net32 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM33<1> net38 net32 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM31 net79 net79 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM4 net_282 PD NEG NEG NHS W=4e-6 L=1e-6 M=1
MM2 PD net4 NEG NEG NHS W=4e-6 L=1e-6 M=1
MM3 PDB PD NEG NEG NHS W=4e-6 L=1e-6 M=1
MM1 net4 PDANA NEG NEG NHS W=4e-6 L=1e-6 M=1
MM73<15> NEG net512 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM73<14> NEG net512 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM73<13> NEG net512 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM73<12> NEG net512 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM73<11> NEG net512 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM73<10> NEG net512 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM73<9> NEG net512 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM73<8> NEG net512 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM73<7> NEG net512 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM73<6> NEG net512 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM73<5> NEG net512 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM73<4> NEG net512 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM73<3> NEG net512 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM73<2> NEG net512 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM73<1> NEG net512 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM73<0> NEG net512 NEG NEG NHS W=4e-6 L=4e-6 M=1
MM5<1> net_282 net512 NEG NEG NHS W=4e-6 L=1e-6 M=1
MM5<0> net_282 net512 NEG NEG NHS W=4e-6 L=1e-6 M=1
MM0 net4 VCOTEST NEG NEG NHS W=4e-6 L=1e-6 M=1
.ENDS

************************************************************************
* Library Name: SINT_mkm18
* Cell Name:    scpllfilt_PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT scpllfilt_PLL600V3_m18 FILPOS FILT FILTER
*.PININFO FILPOS:I FILT:B FILTER:B
RR3 net55 net54 814 $SUB=FILPOS $[R4] $W=2.1e-6 M=1
RR5 net59 net56 814 $SUB=FILPOS $[R4] $W=2.1e-6 M=1
RR2 net54 net49 814 $SUB=FILPOS $[R4] $W=2.1e-6 M=1
RR4 net56 net55 814 $SUB=FILPOS $[R4] $W=2.1e-6 M=1
RR1 net49 net47 814 $SUB=FILPOS $[R4] $W=2.1e-6 M=1
RR7 net1 net61 814 $SUB=FILPOS $[R4] $W=2.1e-6 M=1
RR6 net61 net59 814 $SUB=FILPOS $[R4] $W=2.1e-6 M=1
RR9 FILTER net2 814 $SUB=FILPOS $[R4] $W=2.1e-6 M=1
RR8 net2 net1 814 $SUB=FILPOS $[R4] $W=2.1e-6 M=1
RR0 net47 FILT 814 $SUB=FILPOS $[R4] $W=2.1e-6 M=1
MM1<0> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<1> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<2> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<3> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<4> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<5> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<6> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<7> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<8> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<9> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<10> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<11> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<12> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<13> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<14> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<15> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<16> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<17> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<18> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<19> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<20> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<21> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<22> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<23> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<24> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<25> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<26> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<27> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<28> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<29> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<30> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<31> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<32> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<33> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<34> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<35> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<36> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<37> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<38> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<39> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<40> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<41> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<42> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<43> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<44> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<45> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<46> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<47> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<48> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<49> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<50> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<51> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<52> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<53> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<54> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<55> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<56> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<57> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<58> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<59> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<60> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<61> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<62> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<63> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<64> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<65> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<66> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<67> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<68> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<69> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<70> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<71> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<72> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<73> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<74> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<75> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<76> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<77> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<78> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<79> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<80> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<81> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<82> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<83> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<84> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<85> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<86> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<87> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<88> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<89> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<90> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<91> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<92> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<93> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<94> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<95> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<96> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<97> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<98> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<99> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<100> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<101> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<102> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<103> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<104> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<105> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<106> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<107> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<108> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<109> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<110> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<111> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<112> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<113> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<114> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<115> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<116> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<117> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<118> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<119> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<120> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<121> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<122> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<123> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<124> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<125> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<126> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<127> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<128> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<129> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<130> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<131> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<132> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<133> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<134> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<135> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<136> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<137> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<138> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<139> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<140> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<141> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<142> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<143> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<144> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<145> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<146> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<147> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<148> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<149> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<150> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<151> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<152> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<153> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<154> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<155> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<156> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<157> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<158> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<159> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<160> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<161> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<162> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<163> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<164> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<165> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<166> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<167> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<168> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<169> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<170> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<171> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<172> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<173> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<174> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<175> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<176> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<177> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<178> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<179> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<180> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<181> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<182> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<183> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<184> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<185> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<186> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<187> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<188> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<189> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<190> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<191> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<192> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<193> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<194> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<195> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<196> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<197> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<198> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<199> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<200> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<201> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<202> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<203> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<204> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<205> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<206> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<207> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<208> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<209> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<210> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<211> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<212> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<213> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<214> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<215> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<216> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<217> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<218> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<219> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<220> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<221> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<222> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<223> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<224> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<225> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<226> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<227> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<228> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<229> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<230> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<231> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<232> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<233> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<234> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<235> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<236> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<237> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<238> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<239> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<240> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<241> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<242> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<243> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<244> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<245> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<246> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<247> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<248> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<249> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<250> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<251> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<252> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<253> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<254> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<255> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<256> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<257> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<258> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<259> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<260> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<261> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<262> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<263> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<264> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<265> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<266> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<267> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<268> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<269> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<270> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<271> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<272> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<273> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<274> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<275> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<276> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<277> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<278> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<279> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<280> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<281> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<282> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<283> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<284> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<285> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<286> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<287> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<288> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<289> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<290> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<291> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<292> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<293> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<294> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<295> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<296> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<297> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<298> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<299> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<300> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<301> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<302> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<303> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<304> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<305> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<306> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<307> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<308> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<309> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<310> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<311> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<312> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<313> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<314> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<315> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<316> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<317> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<318> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<319> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<320> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<321> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<322> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<323> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<324> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<325> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<326> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<327> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<328> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<329> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<330> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<331> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<332> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<333> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<334> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<335> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<336> FILPOS FILTER FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM0<0> FILPOS FILT FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM0<1> FILPOS FILT FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM0<2> FILPOS FILT FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM0<3> FILPOS FILT FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM0<4> FILPOS FILT FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM0<5> FILPOS FILT FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM0<6> FILPOS FILT FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM0<7> FILPOS FILT FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM0<8> FILPOS FILT FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM0<9> FILPOS FILT FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
.ENDS

************************************************************************
* Library Name: SINT_mkm18
* Cell Name:    scpllantst_PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT scpllantst_PLL600V3_m18 CHPTEST FREQOK NEG PD POS TESTIO VCOTEST VIN
*.PININFO CHPTEST:I FREQOK:I NEG:I PD:I POS:I VCOTEST:I VIN:I TESTIO:B
XI29 VCOTEST CHPTEST NEG POS net36 / NR2HSP_PLL600V3_m18
MM6 net43 net42 VIN NEG NHS W=0.52e-6 L=0.18e-6 M=1
MM5<0> TESTIO net36 NEG NEG NHS W=1.66e-6 L=0.18e-6 M=1
MM5<1> TESTIO net36 NEG NEG NHS W=1.66e-6 L=0.18e-6 M=1
MM9 VIN net30 TESTIO NEG NHS W=0.52e-6 L=0.18e-6 M=1
MM4<0> net43 net42 TESTIO NEG NHS W=1.66e-6 L=0.18e-6 M=1
MM4<1> net43 net42 TESTIO NEG NHS W=1.66e-6 L=0.18e-6 M=1
MM3<0> TESTIO net85 net43 POS PHS W=1.66e-6 L=0.18e-6 M=1
MM3<1> TESTIO net85 net43 POS PHS W=1.66e-6 L=0.18e-6 M=1
MM7 VIN net85 net43 POS PHS W=0.52e-6 L=0.18e-6 M=1
MM1 VIN FREQOK POS POS PHS W=1.66e-6 L=0.18e-6 M=1
MM8 TESTIO net38 VIN POS PHS W=0.52e-6 L=0.18e-6 M=1
MM0 VIN net78 POS POS PHS W=1.66e-6 L=0.18e-6 M=1
MM2<0> net43 VIN POS POS PHS W=5.74e-6 L=0.5e-6 M=1
MM2<1> net43 VIN POS POS PHS W=5.74e-6 L=0.5e-6 M=1
MM2<2> net43 VIN POS POS PHS W=5.74e-6 L=0.5e-6 M=1
MM2<3> net43 VIN POS POS PHS W=5.74e-6 L=0.5e-6 M=1
MM2<4> net43 VIN POS POS PHS W=5.74e-6 L=0.5e-6 M=1
MM2<5> net43 VIN POS POS PHS W=5.74e-6 L=0.5e-6 M=1
MM2<6> net43 VIN POS POS PHS W=5.74e-6 L=0.5e-6 M=1
MM2<7> net43 VIN POS POS PHS W=5.74e-6 L=0.5e-6 M=1
MM2<8> net43 VIN POS POS PHS W=5.74e-6 L=0.5e-6 M=1
MM2<9> net43 VIN POS POS PHS W=5.74e-6 L=0.5e-6 M=1
MM2<10> net43 VIN POS POS PHS W=5.74e-6 L=0.5e-6 M=1
MM2<11> net43 VIN POS POS PHS W=5.74e-6 L=0.5e-6 M=1
MM2<12> net43 VIN POS POS PHS W=5.74e-6 L=0.5e-6 M=1
MM2<13> net43 VIN POS POS PHS W=5.74e-6 L=0.5e-6 M=1
MM2<14> net43 VIN POS POS PHS W=5.74e-6 L=0.5e-6 M=1
MM2<15> net43 VIN POS POS PHS W=5.74e-6 L=0.5e-6 M=1
XI27 net38 NEG POS net30 / IVHSP_PLL600V3_m18
XI25 VCOTEST NEG POS net85 / IVHSP_PLL600V3_m18
XI26 net85 NEG POS net42 / IVHSP_PLL600V3_m18
XI28 PD NEG POS net78 / IVHSP_PLL600V3_m18
XI24 CHPTEST NEG POS net38 / IVHSP_PLL600V3_m18
.ENDS

************************************************************************
* Library Name: SINT_mkm18
* Cell Name:    DCCV2_2_PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT DCCV2_2_PLL600V3_m18 A NA NEG NY POS Y
*.PININFO A:I NA:I NEG:I POS:I NY:O Y:O
MM6<1> nn2 nn1 NEG NEG NHS W=4e-6 L=0.24e-6 M=1
MM6<0> nn2 nn1 NEG NEG NHS W=4e-6 L=0.24e-6 M=1
MM5<1> n1 n1 NEG NEG NHS W=4e-6 L=0.24e-6 M=1
MM5<0> n1 n1 NEG NEG NHS W=4e-6 L=0.24e-6 M=1
MM12<1> nn1 nn1 NEG NEG NHS W=4e-6 L=0.24e-6 M=1
MM12<0> nn1 nn1 NEG NEG NHS W=4e-6 L=0.24e-6 M=1
MM4<1> n2 n1 NEG NEG NHS W=4e-6 L=0.24e-6 M=1
MM4<0> n2 n1 NEG NEG NHS W=4e-6 L=0.24e-6 M=1
MM3 Y n2 NEG NEG NHS W=1.36e-6 L=0.18e-6 M=1
MM8 NY nn2 NEG NEG NHS W=1.36e-6 L=0.18e-6 M=1
MM11 nn1 A POS POS PHS W=4e-6 L=0.24e-6 M=1
MM1 n2 A POS POS PHS W=4e-6 L=0.24e-6 M=1
MM2 n1 NA POS POS PHS W=4e-6 L=0.24e-6 M=1
MM10 nn2 NA POS POS PHS W=4e-6 L=0.24e-6 M=1
MM9 NY nn2 POS POS PHS W=3.54e-6 L=0.18e-6 M=1
MM0 Y n2 POS POS PHS W=3.54e-6 L=0.18e-6 M=1
.ENDS

************************************************************************
* Library Name: SINT_mkm18
* Cell Name:    PLLVCOMANEATISBIT_2_PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT PLLVCOMANEATISBIT_2_PLL600V3_m18 MINUS NEG OPM OPP PLUS POS Vcn Vcp
*.PININFO MINUS:I NEG:I PLUS:I POS:I Vcn:I Vcp:I OPM:O OPP:O
MM5<1> OPP Vcp POS POS PHS W=6e-6 L=240e-9 M=1
MM5<0> OPP Vcp POS POS PHS W=6e-6 L=240e-9 M=1
MM6 OPP OPP POS POS PHS W=500e-9 L=240e-9 M=1
MM4<1> OPM Vcp POS POS PHS W=6e-6 L=240e-9 M=1
MM4<0> OPM Vcp POS POS PHS W=6e-6 L=240e-9 M=1
MM3 OPM OPM POS POS PHS W=500e-9 L=240e-9 M=1
MM2<1> OPM MINUS net1 NEG NHS W=2.8e-6 L=180e-9 M=1
MM2<0> OPM MINUS net1 NEG NHS W=2.8e-6 L=180e-9 M=1
MM1<1> OPP PLUS net1 NEG NHS W=2.8e-6 L=180e-9 M=1
MM1<0> OPP PLUS net1 NEG NHS W=2.8e-6 L=180e-9 M=1
MM0<3> net1 Vcn NEG NEG NHS W=8e-6 L=240e-9 M=1
MM0<2> net1 Vcn NEG NEG NHS W=8e-6 L=240e-9 M=1
MM0<1> net1 Vcn NEG NEG NHS W=8e-6 L=240e-9 M=1
MM0<0> net1 Vcn NEG NEG NHS W=8e-6 L=240e-9 M=1
.ENDS

************************************************************************
* Library Name: SINT_mkm18
* Cell Name:    PLLVCOMANEATIS_PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT PLLVCOMANEATIS_PLL600V3_m18 CLKR0 NCLKR0 NEG POS Vcp
*.PININFO NEG:I POS:I CLKR0:O NCLKR0:O Vcp:B
DD1 NEG POS DI 1.00e-12
XI58 C0 NC0 NEG NCLKR0 POS CLKR0 / DCCV2_2_PLL600V3_m18
XI62 F<0> NEG NC0 C0 NF<0> POS Vcn Vcp / PLLVCOMANEATISBIT_2_PLL600V3_m18
XI61 F<3> NEG F<0> NF<0> NF<3> POS Vcn Vcp / PLLVCOMANEATISBIT_2_PLL600V3_m18
XI60 F<2> NEG NF<3> F<3> NF<2> POS Vcn Vcp / PLLVCOMANEATISBIT_2_PLL600V3_m18
XI59 F<1> NEG NF<2> F<2> NF<1> POS Vcn Vcp / PLLVCOMANEATISBIT_2_PLL600V3_m18
XI23 F<0> NEG NF<1> F<1> NF<0> POS Vcn Vcp / PLLVCOMANEATISBIT_2_PLL600V3_m18
MM5<3> Vcn Vcn NEG NEG NHS W=8e-6 L=240e-9 M=1
MM5<2> Vcn Vcn NEG NEG NHS W=8e-6 L=240e-9 M=1
MM5<1> Vcn Vcn NEG NEG NHS W=8e-6 L=240e-9 M=1
MM5<0> Vcn Vcn NEG NEG NHS W=8e-6 L=240e-9 M=1
MM4<3> Vcn Vcp POS POS PHS W=6e-6 L=240e-9 M=1
MM4<2> Vcn Vcp POS POS PHS W=6e-6 L=240e-9 M=1
MM4<1> Vcn Vcp POS POS PHS W=6e-6 L=240e-9 M=1
MM4<0> Vcn Vcp POS POS PHS W=6e-6 L=240e-9 M=1
.ENDS

************************************************************************
* Library Name: SERIAL_LINK_mkm18
* Cell Name:    MUX81HSP_PLL600V3_m18
* View Name:    cmos_sch
************************************************************************

.SUBCKT MUX81HSP_PLL600V3_m18 A B C D0 D1 D2 D3 D4 D5 D6 D7 NEG POS Z
*.PININFO A:I B:I C:I D0:I D1:I D2:I D3:I D4:I D5:I D6:I D7:I NEG:I POS:I Z:O
MM144 net1426 net1423 POS POS PHS W=0.62u L=0.18u M=1
MM176 net1419 net2889 net1428 POS PHS W=1.20u L=0.18u M=1
MM140 net2889 net2751 POS POS PHS W=1.24u L=0.18u M=1
MM164 net1431 net2889 net68 POS PHS W=1.20u L=0.18u M=1
MM171 net92 D4 POS POS PHS W=1.20u L=0.18u M=1
MM175 net1428 D6 POS POS PHS W=1.20u L=0.18u M=1
MM168 net1398 net2889 net1316 POS PHS W=1.20u L=0.18u M=1
MM172 net3966 net2889 net92 POS PHS W=1.20u L=0.18u M=1
MM163 net68 D0 POS POS PHS W=1.20u L=0.18u M=1
MM63 net1398 net2751 net86 POS PHS W=1.20u L=0.18u M=1
MM62 net86 D3 POS POS PHS W=1.20u L=0.18u M=1
MM61 net2751 A POS POS PHS W=2.50u L=0.18u M=1
MM60 net1431 net2751 net77 POS PHS W=1.20u L=0.18u M=1
MM59 net77 D1 POS POS PHS W=1.20u L=0.18u M=1
MM181 net3993 net1426 net3966 POS PHS W=1.10u L=0.18u M=1
MM53 Z net120 POS POS PHS W=2.50u L=0.18u M=1
MM52 net118 net1363 POS POS PHS W=0.62u L=0.18u M=1
MM51 net1423 B POS POS PHS W=0.62u L=0.18u M=1
MM50 net120 net1363 net3993 POS PHS W=1.10u L=0.18u M=1
MM48 net3993 net1423 net1419 POS PHS W=1.10u L=0.18u M=1
MM47 net1365 net1423 net1398 POS PHS W=1.10u L=0.18u M=1
MM46 net32 D7 POS POS PHS W=1.20u L=0.18u M=1
MM45 net1419 net2751 net32 POS PHS W=1.20u L=0.18u M=1
MM42 net3966 net2751 net1340 POS PHS W=1.20u L=0.18u M=1
MM41 net1340 D5 POS POS PHS W=1.20u L=0.18u M=1
MM148 net1363 C POS POS PHS W=0.62u L=0.18u M=1
MM167 net1316 D2 POS POS PHS W=1.20u L=0.18u M=1
MM180 net1365 net1426 net1431 POS PHS W=1.10u L=0.18u M=1
MM183 net120 net118 net1365 POS PHS W=1.10u L=0.18u M=1
MM166 net1434 D0 NEG NEG NHS W=0.52u L=0.18u M=1
MM165 net1431 net2751 net1434 NEG NHS W=0.52u L=0.18u M=1
MM87 net1422 D7 NEG NEG NHS W=0.52u L=0.18u M=1
MM86 net1419 net2889 net1422 NEG NHS W=0.52u L=0.18u M=1
MM83 net1410 D5 NEG NEG NHS W=0.52u L=0.18u M=1
MM82 net3966 net2889 net1410 NEG NHS W=0.52u L=0.18u M=1
MM79 net1398 net2889 net1395 NEG NHS W=0.52u L=0.18u M=1
MM77 net2751 A NEG NEG NHS W=1.42u L=0.18u M=1
MM76 net1392 D1 NEG NEG NHS W=0.52u L=0.18u M=1
MM75 net1431 net2889 net1392 NEG NHS W=0.52u L=0.18u M=1
MM71 Z net120 NEG NEG NHS W=1.42u L=0.18u M=1
MM70 net118 net1363 NEG NEG NHS W=0.34u L=0.18u M=1
MM69 net1423 B NEG NEG NHS W=0.34u L=0.18u M=1
MM68 net120 net118 net3993 NEG NHS W=0.84u L=0.20u M=1
MM66 net1365 net1426 net1398 NEG NHS W=0.84u L=0.20u M=1
MM174 net1404 D4 NEG NEG NHS W=0.52u L=0.18u M=1
MM173 net3966 net2751 net1404 NEG NHS W=0.52u L=0.18u M=1
MM169 net1398 net2751 net1383 NEG NHS W=0.52u L=0.18u M=1
MM177 net1419 net2751 net1416 NEG NHS W=0.52u L=0.18u M=1
MM178 net1416 D6 NEG NEG NHS W=0.52u L=0.18u M=1
MM170 net1383 D2 NEG NEG NHS W=0.52u L=0.18u M=1
MM141 net2889 net2751 NEG NEG NHS W=0.70u L=0.18u M=1
MM145 net1426 net1423 NEG NEG NHS W=0.34u L=0.18u M=1
MM149 net1363 C NEG NEG NHS W=0.34u L=0.18u M=1
MM156 net1395 D3 NEG NEG NHS W=0.52u L=0.18u M=1
MM184 net120 net1363 net1365 NEG NHS W=0.84u L=0.20u M=1
MM182 net3993 net1423 net3966 NEG NHS W=0.84u L=0.20u M=1
MM179 net1365 net1423 net1431 NEG NHS W=0.84u L=0.20u M=1
MM89 net3993 net1426 net1419 NEG NHS W=0.84u L=0.20u M=1
DD227 A POS DP 1.02e-13
DD189 D6 POS DP 1.02e-13
DD221 NEG D0 DN 1.02e-13
DD217 NEG D1 DN 1.02e-13
DD213 NEG C DN 1.02e-13
DD209 NEG B DN 1.02e-13
DD205 NEG D2 DN 1.02e-13
DD201 NEG D3 DN 1.02e-13
DD197 NEG D4 DN 1.02e-13
DD193 NEG D5 DN 1.02e-13
DD185 NEG D7 DN 1.02e-13
.ENDS

************************************************************************
* Library Name: SINT_mkm18
* Cell Name:    scpllopdvb_PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT scpllopdvb_PLL600V3_m18 CLK CLKB NEG POS Q QB TOG
*.PININFO CLK:I CLKB:I NEG:I POS:I TOG:I Q:O QB:O
MM14 net165 net162 POS POS PHS W=1.66e-6 L=0.18e-6 M=1
MM13 Q QB POS POS PHS W=1.66e-6 L=0.18e-6 M=1
MM29 QB Q POS POS PHS W=1.66e-6 L=0.18e-6 M=1
MM30 net162 net165 POS POS PHS W=1.66e-6 L=0.18e-6 M=1
MM12 net165 net162 NEG NEG NHS W=0.52e-6 L=0.18e-6 M=1
MM33 QB CLK net48 NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM25 net120 Q net117 NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM9 net96 TOG NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM7 net99 QB net96 NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM8 net36 QB net89 NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM21 net86 TOG NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM38 net87 net162 NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM34 QB CLK net108 NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM32 net108 net165 NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM10 net89 TOG NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM22 net39 Q net86 NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM11 Q QB NEG NEG NHS W=0.52e-6 L=0.18e-6 M=1
MM6 net162 CLKB net36 NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM23 net165 CLKB net39 NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM36 Q CLK net51 NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM35 Q CLK net87 NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM28 net162 net165 NEG NEG NHS W=0.52e-6 L=0.18e-6 M=1
MM37 net51 net162 NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM27 QB Q NEG NEG NHS W=0.52e-6 L=0.18e-6 M=1
MM5 net162 CLKB net99 NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM24 net117 TOG NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM31 net48 net165 NEG NEG NHS W=1.56e-6 L=0.18e-6 M=1
MM26 net165 CLKB net120 NEG NHS W=1.56e-6 L=0.18e-6 M=1
.ENDS

************************************************************************
* Library Name: SINT_mkm18
* Cell Name:    scpllopdiv_PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT scpllopdiv_PLL600V3_m18 BYPASS CLKBYP CLKIN CLKOUTB DV0 DV1 FORCE1 NEG 
+ POS
*.PININFO BYPASS:I CLKBYP:I CLKIN:I DV0:I DV1:I FORCE1:I NEG:I POS:I CLKOUTB:O
XI61 net1 net4 net2 NEG POS Y2 / AN3HSP_PLL600V3_m18
XI60 net1 net3 net2 NEG POS Y1 / AN3HSP_PLL600V3_m18
XI48 Y1 Y2 Y3 CLKIN divide2 divide4 divide8 net154 TIELO TIELO TIELO NEG POS 
+ net5 / MUX81HSP_PLL600V3_m18
XI36 NEG POS TIELO / TIELO_PLL600V3_m18
XI23 CLK CLKB NEG POS net122 net13 divide2 / scpllopdvb_PLL600V3_m18
XI24 CLK CLKB NEG POS net116 net7 net394 / scpllopdvb_PLL600V3_m18
XXI1 CLK CLKB NEG POS net128 net25 POS / scpllopdvb_PLL600V3_m18
XI21 net128 net122 NEG POS net394 / AN2HSP_PLL600V3_m18
XI18 CLKBYP NEG POS net154 / IVHSX4_PLL600V3_m18
XI58 net5 NEG POS CLKOUTB / IVHSX4_PLL600V3_m18
XI9 net13 NEG POS divide4 / IVHSP_PLL600V3_m18
XI8 net25 NEG POS divide2 / IVHSP_PLL600V3_m18
XI12 net7 NEG POS divide8 / IVHSP_PLL600V3_m18
XI53 DV0 NEG POS net8 / IVHSP_PLL600V3_m18
XI64 net8 NEG POS net3 / IVHSP_PLL600V3_m18
XI54 FORCE1 NEG POS net1 / IVHSP_PLL600V3_m18
XI50 BYPASS NEG POS net2 / IVHSP_PLL600V3_m18
XI63 net6 NEG POS net4 / IVHSP_PLL600V3_m18
XI7 CLKIN NEG POS CLKB / IVHSP_PLL600V3_m18
XI6 net343 NEG POS CLK / IVHSP_PLL600V3_m18
XI5 CLKIN NEG POS net343 / IVHSP_PLL600V3_m18
XI51 DV1 NEG POS net6 / IVHSP_PLL600V3_m18
XI62 net2 NEG POS Y3 / IVHSP_PLL600V3_m18
.ENDS

************************************************************************
* Library Name: SERIAL_LINK_mkm18
* Cell Name:    MXI2HSX2_PLL600V3_m18
* View Name:    cmos_sch
************************************************************************

.SUBCKT MXI2HSX2_PLL600V3_m18 A B NEG POS S0 Y
*.PININFO A:I B:I NEG:I POS:I S0:I Y:O
MMN3 net3 B NEG NEG NHS W=1.56u L=0.18u M=1
MMN4 Y S0 net3 NEG NHS W=1.56u L=0.18u M=1
MMN2 Y net660 net12 NEG NHS W=1.56u L=0.18u M=1
MMN1 net12 A NEG NEG NHS W=1.56u L=0.18u M=1
MMN29 net660 S0 NEG NEG NHS W=1.14u L=0.18u M=1
MMP4 Y net660 net622 POS PHS W=2.20u L=0.18u M=1
MMP3 Y S0 net18 POS PHS W=2.20u L=0.18u M=1
MMP2 net622 B POS POS PHS W=2.20u L=0.18u M=1
MMP1 net18 A POS POS PHS W=2.20u L=0.18u M=1
MMP28 net660 S0 POS POS PHS W=1.46u L=0.18u M=1
DD32 B POS DP 1.02e-13
DD0 A POS DP 1.02e-13
DD40 NEG S0 DN 1.02e-13
.ENDS

************************************************************************
* Library Name: SINT_mkm18
* Cell Name:    pllfcs_fix1_PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT pllfcs_fix1_PLL600V3_m18 BYPASS CLKBYP CLKCONTR CLKCORE CLKDDRIN 
+ CLKDDROUT CLKIN FORCE1 NEG POS SLOW_MEM
*.PININFO BYPASS:I CLKBYP:I CLKIN:I FORCE1:I NEG:I POS:I SLOW_MEM:I CLKCONTR:O 
*.PININFO CLKCORE:O CLKDDRIN:O CLKDDROUT:O
XI270 NEG POS TIELO / TIELO_PLL600V3_m18
XI254 net0111 net0106 NEG POS net096 / ND2HSP_PLL600V3_m18
XI250 net0270 net0120 NEG POS net0105 / ND2HSP_PLL600V3_m18
XI248 net0118 net0113 NEG POS net0107 / ND2HSP_PLL600V3_m18
XI253 net0105 net0121 NEG POS net0106 / ND2HSP_PLL600V3_m18
XI252 net0110 net0263 NEG POS net0111 / ND2HSP_PLL600V3_m18
XI246 net089 net0270 NEG POS net0118 / ND2HSP_PLL600V3_m18
XI247 net0286 net0120 NEG POS net0113 / ND2HSP_PLL600V3_m18
XI249 net0270 net0120 NEG POS net0179 net0133 S / FD4HSP_PLL600V3_m18
XI257 CLK net096 NEG POS net0104 net0176 S / FD4HSP_PLL600V3_m18
XI268 CLK net4 NEG POS CLKCONTR net5 S / FD4HSP_PLL600V3_m18
XI258 net0260 net0121 NEG POS net0156 net0188 S / FD4HSP_PLL600V3_m18
XI267 CLK net2 NEG POS CLKDDROUT net3 S / FD4HSP_PLL600V3_m18
XI245 CLK net0107 NEG POS net0260 net0139 S / FD4HSP_PLL600V3_m18
XI244 CLK net0190 NEG POS net087 net0192 S / FD4HSP_PLL600V3_m18
XI266 CLK net0247 NEG POS CLKCORE net1 S / FD4HSP_PLL600V3_m18
XI269 CLK net080 NEG POS CLKDDRIN net058 S / FD4HSP_PLL600V3_m18
XI241 net0179 NEG POS net095 / IVHSP_PLL600V3_m18
XI238 net0260 NEG POS net089 / IVHSP_PLL600V3_m18
XI240 net0139 NEG POS net0120 / IVHSP_PLL600V3_m18
XI235 net087 NEG POS net0270 / IVHSP_PLL600V3_m18
XI255 net0104 NEG POS net0110 / IVHSP_PLL600V3_m18
XI256 net0176 NEG POS net0121 / IVHSP_PLL600V3_m18
XI251 net0105 NEG POS net0263 / IVHSP_PLL600V3_m18
XI239 net0260 NEG POS net0257 / IVHSP_PLL600V3_m18
XI233 net0100 NEG POS CLK / IVHSP_PLL600V3_m18
XI236 net0192 NEG POS net0286 / IVHSP_PLL600V3_m18
XI234 net087 NEG POS net0190 / IVHSP_PLL600V3_m18
XI237 FORCE1 NEG POS S / IVHSX4_PLL600V3_m18
XI231 net0112 NEG POS net0318 / IVHSX4_PLL600V3_m18
XI271 SLOW_MEM NEG POS net0108 / IVHSX4_PLL600V3_m18
XI272 net0108 NEG POS net6 / IVHSX4_PLL600V3_m18
XI230 BYPASS NEG POS net0112 / IVHSX4_PLL600V3_m18
XI284 net0286 TIELO NEG POS TIELO net0247 / MXI2HSX2_PLL600V3_m18
XI287 net095 net0156 NEG POS net6 net080 / MXI2HSX2_PLL600V3_m18
XI285 net0286 net0257 NEG POS net6 net2 / MXI2HSX2_PLL600V3_m18
XI290 CLKIN CLKBYP NEG POS net0318 net0100 / MXI2HSX2_PLL600V3_m18
XI286 net0257 net0121 NEG POS net6 net4 / MXI2HSX2_PLL600V3_m18
.ENDS

************************************************************************
* Library Name: SINT_mkm18
* Cell Name:    PLL600V3_m18
* View Name:    schematic
************************************************************************

.SUBCKT PLL600V3_m18 AT1 BMCLK1X CHP0 CHP1 CHP2 CHP3 CHP4 
+ CLKCONTR CLKCORE CLKDDRIN CLKDDROUT CLKFBKB DIV0 DIV1 DIV2 DIV3 DIV4 DT1 ENB 
+ LKDET PD PLLGND PLLVDD SG1 SLOW_MEM SYNCEN TM1 TM2 VCOD0 VCOD1
*.PININFO BMCLK1X:I CHP0:I CHP1:I CHP2:I CHP3:I CHP4:I CLKFBKB:I DIV0:I DIV1:I 
*.PININFO DIV2:I DIV3:I DIV4:I ENB:I PD:I SG1:I SLOW_MEM:I SYNCEN:I TM1:I 
*.PININFO TM2:I VCOD0:I VCOD1:I AT1:O CLKCONTR:O CLKCORE:O CLKDDRIN:O 
*.PININFO CLKDDROUT:O DT1:O LKDET:O PLLGND:B PLLVDD:B
XI81 C2 CLKFDB2 IBIAS PLLGND PDANA PLLVDD TM1 / scpllochk_V2_PLL600V3_m18
XI120 net0119 PLLGND PLLVDD CLKDDRIN / IVHSP_PLL600V3_m18
XI119 net0121 PLLGND PLLVDD CLKCONTR / IVHSP_PLL600V3_m18
XI118 net0122 PLLGND PLLVDD CLKDDROUT / IVHSP_PLL600V3_m18
XI117 net0120 PLLGND PLLVDD CLKCORE / IVHSP_PLL600V3_m18
XI111 net0128 PLLGND PLLVDD BNMCLK1X / IVHSP_PLL600V3_m18
XI109 net0129 PLLGND PLLVDD CLKFDB2 / IVHSP_PLL600V3_m18
XI110 net098 PLLGND PLLVDD net0128 / IVHSP_PLL600V3_m18
XI108 net097 PLLGND PLLVDD net0129 / IVHSP_PLL600V3_m18
XI114 BMCLK1X PLLGND PLLVDD net098 / IVHSP_PLL600V3_m18
XI115 CLKFBKB PLLGND PLLVDD net097 / IVHSP_PLL600V3_m18
XI83 net097 DIV0 DIV1 DIV2 DIV3 DIV4 CLKFDB net073 FORCE32 PLLGND PLLVDD 
+ DIVRES SYNCEN / scplldivid_PLL600V3_m18
XI82 net098 PLLGND PLLGND PLLGND PLLGND PLLGND net0109 net0132 PLLGND PLLGND 
+ PLLVDD DIVRES PLLVDD / scplldivid_PLL600V3_m18
XI123 FILPOS PLLGND PLLVDD / PLLFILTSUPV2_PLL600V3_m18
XI95 CLKBCKB CLKFDB net0109 CLKREFB PLLGND PLLVDD CHPTEST SG1 / 
+ pllipmux_PLL600V3_m18
XI85 BNMCLK1X INTDT1 PLLGND DT1 PLLVDD SG1 TM1 TM2 / scplltfac_PLL600V3_m18
XI79 CHPTEST net073 DIVRES INTDT1 ENB FORCE32 PLLGND PD PDANA PLLVDD SG1 TM1 
+ TM2 VCOTEST / scplltcon_PLL600V3_m18
XI76 CLKBCKB CLKREFB DN DNB net0125 net0126 PLLGND net0123 net0124 PLLVDD UP 
+ UPB / scpllphdet_PLL600V3_m18
MM1<0> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<1> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<2> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<3> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<4> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<5> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<6> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<7> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<8> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<9> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<10> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<11> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<12> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<13> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<14> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<15> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<16> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<17> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<18> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<19> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<20> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<21> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<22> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<23> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<24> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<25> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<26> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<27> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<28> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<29> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<30> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<31> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<32> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<33> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<34> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<35> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<36> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<37> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<38> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<39> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<40> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<41> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<42> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<43> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<44> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<45> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<46> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<47> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<48> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<49> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<50> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<51> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<52> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<53> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<54> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<55> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<56> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<57> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<58> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<59> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<60> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<61> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<62> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<63> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<64> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<65> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<66> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<67> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<68> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<69> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<70> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<71> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<72> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<73> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<74> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<75> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<76> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<77> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<78> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<79> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<80> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<81> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<82> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<83> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<84> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<85> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<86> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<87> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<88> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<89> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<90> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<91> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<92> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<93> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<94> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<95> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<96> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<97> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<98> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<99> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<100> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<101> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<102> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<103> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<104> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<105> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<106> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<107> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<108> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<109> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<110> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<111> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<112> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<113> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<114> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<115> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<116> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM1<117> FILPOS PLLGND FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<0> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<1> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<2> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<3> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<4> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<5> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<6> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<7> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<8> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<9> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<10> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<11> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<12> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<13> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<14> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<15> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<16> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<17> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<18> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<19> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<20> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<21> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<22> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<23> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<24> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<25> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<26> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<27> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<28> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<29> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<30> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<31> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<32> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<33> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<34> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<35> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<36> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<37> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<38> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<39> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<40> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<41> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<42> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<43> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<44> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<45> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<46> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<47> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<48> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<49> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<50> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<51> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<52> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<53> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<54> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<55> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<56> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<57> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<58> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<59> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<60> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<61> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<62> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<63> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<64> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<65> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<66> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<67> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<68> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<69> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<70> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<71> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<72> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<73> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<74> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<75> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<76> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<77> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<78> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<79> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<80> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<81> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<82> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<83> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<84> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<85> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<86> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<87> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<88> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<89> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<90> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<91> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<92> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<93> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<94> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<95> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<96> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<97> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<98> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<99> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<100> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<101> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<102> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<103> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<104> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
MM2<105> FILPOS net0131 FILPOS FILPOS PHS W=9.4e-6 L=4.54e-6 M=1
XI107 LKDET net0125 net0126 PLLGND PDANA net0123 net0124 PLLVDD / 
+ scplllkdet_PLL600V3_m18
XI78 net0131 CHP0 CHP1 CHP2 CHP3 CHP4 VIN DN DNB IBIAS PLLGND PDANA FILPOS UP 
+ UPB VCOTEST / scpllchgpmp_PLL600V3_m18
XI86 FILPOS VIN C2 / scpllfilt_PLL600V3_m18
XI77 CHPTEST PLLVDD PLLGND PDANA FILPOS AT1 VCOTEST VIN / 
+ scpllantst_PLL600V3_m18
DD0 PLLGND FILPOS DI 1.00e-12
DD1 PLLGND PLLVDD DI 1.00e-12
XI121 VCOOUT net0133 PLLGND FILPOS VIN / PLLVCOMANEATIS_PLL600V3_m18
XI101 PLLGND PLLGND VCOOUT net0118 VCOD0 VCOD1 PDANA PLLGND PLLVDD / 
+ scpllopdiv_PLL600V3_m18
XI87 TM2 BNMCLK1X net0121 net0120 net0119 net0122 net0118 PD PLLGND PLLVDD 
+ SLOW_MEM / pllfcs_fix1_PLL600V3_m18
.ENDS

