//--------------------------------------------------------------------------------
// 
//              Verilog models for the CORELIB8DHS.HCMOS8D
//                    (CORELIB8DHS)
// 
//
//--------------------------------------------------------------------------------
// CELL AN2HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN2HS_B_F_Z_F 0.1
`define AN2HS_B_R_Z_R 0.1
`define AN2HS_A_F_Z_F 0.1
`define AN2HS_A_R_Z_R 0.1

module AN2HS (Z, A, B);

   output Z;
   input A;
   input B;


   and  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B +=> Z) = (`AN2HS_B_R_Z_R,`AN2HS_B_F_Z_F);
      (A +=> Z) = (`AN2HS_A_R_Z_R,`AN2HS_A_F_Z_F);

   endspecify
`endif


endmodule // AN2HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:46 and Version :1.1 //
 
//  START 
// CELL AN2HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN2HSP_B_F_Z_F 0.1
`define AN2HSP_B_R_Z_R 0.1
`define AN2HSP_A_F_Z_F 0.1
`define AN2HSP_A_R_Z_R 0.1

module AN2HSP (Z, A, B);

   output Z;
   input A;
   input B;


   and  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B +=> Z) = (`AN2HSP_B_R_Z_R,`AN2HSP_B_F_Z_F);
      (A +=> Z) = (`AN2HSP_A_R_Z_R,`AN2HSP_A_F_Z_F);

   endspecify
`endif


endmodule // AN2HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:46 and Version :1.1 //
 
//  START 
// CELL AN2HSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN2HSX3_B_F_Z_F 0.1
`define AN2HSX3_B_R_Z_R 0.1
`define AN2HSX3_A_F_Z_F 0.1
`define AN2HSX3_A_R_Z_R 0.1

module AN2HSX3 (Z, A, B);

   output Z;
   input A;
   input B;


   and  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B +=> Z) = (`AN2HSX3_B_R_Z_R,`AN2HSX3_B_F_Z_F);
      (A +=> Z) = (`AN2HSX3_A_R_Z_R,`AN2HSX3_A_F_Z_F);

   endspecify
`endif


endmodule // AN2HSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:46 and Version :1.1 //
 
//  START 
// CELL AN2HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN2HSX4_B_F_Z_F 0.1
`define AN2HSX4_B_R_Z_R 0.1
`define AN2HSX4_A_F_Z_F 0.1
`define AN2HSX4_A_R_Z_R 0.1

module AN2HSX4 (Z, A, B);

   output Z;
   input A;
   input B;


   and  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B +=> Z) = (`AN2HSX4_B_R_Z_R,`AN2HSX4_B_F_Z_F);
      (A +=> Z) = (`AN2HSX4_A_R_Z_R,`AN2HSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AN2HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:46 and Version :1.1 //
 
//  START 
// CELL AN2HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN2HSX8_B_F_Z_F 0.1
`define AN2HSX8_B_R_Z_R 0.1
`define AN2HSX8_A_F_Z_F 0.1
`define AN2HSX8_A_R_Z_R 0.1

module AN2HSX8 (Z, A, B);

   output Z;
   input A;
   input B;


   and  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B +=> Z) = (`AN2HSX8_B_R_Z_R,`AN2HSX8_B_F_Z_F);
      (A +=> Z) = (`AN2HSX8_A_R_Z_R,`AN2HSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AN2HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:46 and Version :1.1 //
 
//  START 
// CELL F_AN2HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AN2HSP_B_F_Z_F 0.1
`define F_AN2HSP_B_R_Z_R 0.1
`define F_AN2HSP_A_F_Z_F 0.1
`define F_AN2HSP_A_R_Z_R 0.1

module F_AN2HSP (Z, A, B);

   output Z;
   input A;
   input B;


   and  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B +=> Z) = (`F_AN2HSP_B_R_Z_R,`F_AN2HSP_B_F_Z_F);
      (A +=> Z) = (`F_AN2HSP_A_R_Z_R,`F_AN2HSP_A_F_Z_F);

   endspecify
`endif


endmodule // F_AN2HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:46 and Version :1.1 //
 
//  START 
// CELL AN2AHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN2AHS_B_F_Z_F 0.1
`define AN2AHS_B_R_Z_R 0.1
`define AN2AHS_A_F_Z_R 0.1
`define AN2AHS_A_R_Z_F 0.1

module AN2AHS (Z, A, B);

   output Z;
   input A;
   input B;


   and  u0 (Z, AX, B);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (B +=> Z) = (`AN2AHS_B_R_Z_R,`AN2AHS_B_F_Z_F);
      (A -=> Z) = (`AN2AHS_A_F_Z_R,`AN2AHS_A_R_Z_F);

   endspecify
`endif


endmodule // AN2AHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:46 and Version :1.1 //
 
//  START 
// CELL AN2AHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN2AHSP_B_F_Z_F 0.1
`define AN2AHSP_B_R_Z_R 0.1
`define AN2AHSP_A_F_Z_R 0.1
`define AN2AHSP_A_R_Z_F 0.1

module AN2AHSP (Z, A, B);

   output Z;
   input A;
   input B;


   and  u0 (Z, AX, B);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (B +=> Z) = (`AN2AHSP_B_R_Z_R,`AN2AHSP_B_F_Z_F);
      (A -=> Z) = (`AN2AHSP_A_F_Z_R,`AN2AHSP_A_R_Z_F);

   endspecify
`endif


endmodule // AN2AHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:46 and Version :1.1 //
 
//  START 
// CELL AN2AHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN2AHSX4_B_F_Z_F 0.1
`define AN2AHSX4_B_R_Z_R 0.1
`define AN2AHSX4_A_F_Z_R 0.1
`define AN2AHSX4_A_R_Z_F 0.1

module AN2AHSX4 (Z, A, B);

   output Z;
   input A;
   input B;


   and  u0 (Z, AX, B);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (B +=> Z) = (`AN2AHSX4_B_R_Z_R,`AN2AHSX4_B_F_Z_F);
      (A -=> Z) = (`AN2AHSX4_A_F_Z_R,`AN2AHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AN2AHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:46 and Version :1.1 //
 
//  START 
// CELL AN3HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN3HS_C_F_Z_F 0.1
`define AN3HS_C_R_Z_R 0.1
`define AN3HS_B_F_Z_F 0.1
`define AN3HS_B_R_Z_R 0.1
`define AN3HS_A_F_Z_F 0.1
`define AN3HS_A_R_Z_R 0.1

module AN3HS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AN3HS_C_R_Z_R,`AN3HS_C_F_Z_F);
      (B +=> Z) = (`AN3HS_B_R_Z_R,`AN3HS_B_F_Z_F);
      (A +=> Z) = (`AN3HS_A_R_Z_R,`AN3HS_A_F_Z_F);

   endspecify
`endif


endmodule // AN3HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:51 and Version :1.1 //
 
//  START 
// CELL AN3HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN3HSP_C_F_Z_F 0.1
`define AN3HSP_C_R_Z_R 0.1
`define AN3HSP_B_F_Z_F 0.1
`define AN3HSP_B_R_Z_R 0.1
`define AN3HSP_A_F_Z_F 0.1
`define AN3HSP_A_R_Z_R 0.1

module AN3HSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AN3HSP_C_R_Z_R,`AN3HSP_C_F_Z_F);
      (B +=> Z) = (`AN3HSP_B_R_Z_R,`AN3HSP_B_F_Z_F);
      (A +=> Z) = (`AN3HSP_A_R_Z_R,`AN3HSP_A_F_Z_F);

   endspecify
`endif


endmodule // AN3HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:51 and Version :1.1 //
 
//  START 
// CELL AN3HSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN3HSX3_C_F_Z_F 0.1
`define AN3HSX3_C_R_Z_R 0.1
`define AN3HSX3_B_F_Z_F 0.1
`define AN3HSX3_B_R_Z_R 0.1
`define AN3HSX3_A_F_Z_F 0.1
`define AN3HSX3_A_R_Z_R 0.1

module AN3HSX3 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AN3HSX3_C_R_Z_R,`AN3HSX3_C_F_Z_F);
      (B +=> Z) = (`AN3HSX3_B_R_Z_R,`AN3HSX3_B_F_Z_F);
      (A +=> Z) = (`AN3HSX3_A_R_Z_R,`AN3HSX3_A_F_Z_F);

   endspecify
`endif


endmodule // AN3HSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:51 and Version :1.1 //
 
//  START 
// CELL AN3HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN3HSX4_C_F_Z_F 0.1
`define AN3HSX4_C_R_Z_R 0.1
`define AN3HSX4_B_F_Z_F 0.1
`define AN3HSX4_B_R_Z_R 0.1
`define AN3HSX4_A_F_Z_F 0.1
`define AN3HSX4_A_R_Z_R 0.1

module AN3HSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AN3HSX4_C_R_Z_R,`AN3HSX4_C_F_Z_F);
      (B +=> Z) = (`AN3HSX4_B_R_Z_R,`AN3HSX4_B_F_Z_F);
      (A +=> Z) = (`AN3HSX4_A_R_Z_R,`AN3HSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AN3HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:51 and Version :1.1 //
 
//  START 
// CELL AN3HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN3HSX8_C_F_Z_F 0.1
`define AN3HSX8_C_R_Z_R 0.1
`define AN3HSX8_B_F_Z_F 0.1
`define AN3HSX8_B_R_Z_R 0.1
`define AN3HSX8_A_F_Z_F 0.1
`define AN3HSX8_A_R_Z_R 0.1

module AN3HSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AN3HSX8_C_R_Z_R,`AN3HSX8_C_F_Z_F);
      (B +=> Z) = (`AN3HSX8_B_R_Z_R,`AN3HSX8_B_F_Z_F);
      (A +=> Z) = (`AN3HSX8_A_R_Z_R,`AN3HSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AN3HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:51 and Version :1.1 //
 
//  START 
// CELL AN3AHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN3AHS_C_F_Z_F 0.1
`define AN3AHS_C_R_Z_R 0.1
`define AN3AHS_B_F_Z_F 0.1
`define AN3AHS_B_R_Z_R 0.1
`define AN3AHS_A_F_Z_R 0.1
`define AN3AHS_A_R_Z_F 0.1

module AN3AHS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AN3AHS_C_R_Z_R,`AN3AHS_C_F_Z_F);
      (B +=> Z) = (`AN3AHS_B_R_Z_R,`AN3AHS_B_F_Z_F);
      (A -=> Z) = (`AN3AHS_A_F_Z_R,`AN3AHS_A_R_Z_F);

   endspecify
`endif


endmodule // AN3AHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:51 and Version :1.1 //
 
//  START 
// CELL AN3AHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN3AHSP_C_F_Z_F 0.1
`define AN3AHSP_C_R_Z_R 0.1
`define AN3AHSP_B_F_Z_F 0.1
`define AN3AHSP_B_R_Z_R 0.1
`define AN3AHSP_A_F_Z_R 0.1
`define AN3AHSP_A_R_Z_F 0.1

module AN3AHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AN3AHSP_C_R_Z_R,`AN3AHSP_C_F_Z_F);
      (B +=> Z) = (`AN3AHSP_B_R_Z_R,`AN3AHSP_B_F_Z_F);
      (A -=> Z) = (`AN3AHSP_A_F_Z_R,`AN3AHSP_A_R_Z_F);

   endspecify
`endif


endmodule // AN3AHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:51 and Version :1.1 //
 
//  START 
// CELL AN3AHSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN3AHSX3_C_F_Z_F 0.1
`define AN3AHSX3_C_R_Z_R 0.1
`define AN3AHSX3_B_F_Z_F 0.1
`define AN3AHSX3_B_R_Z_R 0.1
`define AN3AHSX3_A_F_Z_R 0.1
`define AN3AHSX3_A_R_Z_F 0.1

module AN3AHSX3 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AN3AHSX3_C_R_Z_R,`AN3AHSX3_C_F_Z_F);
      (B +=> Z) = (`AN3AHSX3_B_R_Z_R,`AN3AHSX3_B_F_Z_F);
      (A -=> Z) = (`AN3AHSX3_A_F_Z_R,`AN3AHSX3_A_R_Z_F);

   endspecify
`endif


endmodule // AN3AHSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:51 and Version :1.1 //
 
//  START 
// CELL AN3AHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN3AHSX4_C_F_Z_F 0.1
`define AN3AHSX4_C_R_Z_R 0.1
`define AN3AHSX4_B_F_Z_F 0.1
`define AN3AHSX4_B_R_Z_R 0.1
`define AN3AHSX4_A_F_Z_R 0.1
`define AN3AHSX4_A_R_Z_F 0.1

module AN3AHSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AN3AHSX4_C_R_Z_R,`AN3AHSX4_C_F_Z_F);
      (B +=> Z) = (`AN3AHSX4_B_R_Z_R,`AN3AHSX4_B_F_Z_F);
      (A -=> Z) = (`AN3AHSX4_A_F_Z_R,`AN3AHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AN3AHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:51 and Version :1.1 //
 
//  START 
// CELL AN3AHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN3AHSX8_C_F_Z_F 0.1
`define AN3AHSX8_C_R_Z_R 0.1
`define AN3AHSX8_B_F_Z_F 0.1
`define AN3AHSX8_B_R_Z_R 0.1
`define AN3AHSX8_A_F_Z_R 0.1
`define AN3AHSX8_A_R_Z_F 0.1

module AN3AHSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AN3AHSX8_C_R_Z_R,`AN3AHSX8_C_F_Z_F);
      (B +=> Z) = (`AN3AHSX8_B_R_Z_R,`AN3AHSX8_B_F_Z_F);
      (A -=> Z) = (`AN3AHSX8_A_F_Z_R,`AN3AHSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AN3AHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:51 and Version :1.1 //
 
//  START 
// CELL AN4HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN4HS_D_F_Z_F 0.1
`define AN4HS_D_R_Z_R 0.1
`define AN4HS_C_F_Z_F 0.1
`define AN4HS_C_R_Z_R 0.1
`define AN4HS_B_F_Z_F 0.1
`define AN4HS_B_R_Z_R 0.1
`define AN4HS_A_F_Z_F 0.1
`define AN4HS_A_R_Z_R 0.1

module AN4HS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AN4HS_D_R_Z_R,`AN4HS_D_F_Z_F);
      (C +=> Z) = (`AN4HS_C_R_Z_R,`AN4HS_C_F_Z_F);
      (B +=> Z) = (`AN4HS_B_R_Z_R,`AN4HS_B_F_Z_F);
      (A +=> Z) = (`AN4HS_A_R_Z_R,`AN4HS_A_F_Z_F);

   endspecify
`endif


endmodule // AN4HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:54 and Version :1.1 //

//  START
// CELL AN4HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN4HSP_D_F_Z_F 0.1
`define AN4HSP_D_R_Z_R 0.1
`define AN4HSP_C_F_Z_F 0.1
`define AN4HSP_C_R_Z_R 0.1
`define AN4HSP_B_F_Z_F 0.1
`define AN4HSP_B_R_Z_R 0.1
`define AN4HSP_A_F_Z_F 0.1
`define AN4HSP_A_R_Z_R 0.1

module AN4HSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AN4HSP_D_R_Z_R,`AN4HSP_D_F_Z_F);
      (C +=> Z) = (`AN4HSP_C_R_Z_R,`AN4HSP_C_F_Z_F);
      (B +=> Z) = (`AN4HSP_B_R_Z_R,`AN4HSP_B_F_Z_F);
      (A +=> Z) = (`AN4HSP_A_R_Z_R,`AN4HSP_A_F_Z_F);

   endspecify
`endif


endmodule // AN4HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:54 and Version :1.1 //

//  START
// CELL AN4HSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN4HSX3_D_F_Z_F 0.1
`define AN4HSX3_D_R_Z_R 0.1
`define AN4HSX3_C_F_Z_F 0.1
`define AN4HSX3_C_R_Z_R 0.1
`define AN4HSX3_B_F_Z_F 0.1
`define AN4HSX3_B_R_Z_R 0.1
`define AN4HSX3_A_F_Z_F 0.1
`define AN4HSX3_A_R_Z_R 0.1

module AN4HSX3 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AN4HSX3_D_R_Z_R,`AN4HSX3_D_F_Z_F);
      (C +=> Z) = (`AN4HSX3_C_R_Z_R,`AN4HSX3_C_F_Z_F);
      (B +=> Z) = (`AN4HSX3_B_R_Z_R,`AN4HSX3_B_F_Z_F);
      (A +=> Z) = (`AN4HSX3_A_R_Z_R,`AN4HSX3_A_F_Z_F);

   endspecify
`endif


endmodule // AN4HSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:54 and Version :1.1 //

//  START
// CELL AN4HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN4HSX4_D_F_Z_F 0.1
`define AN4HSX4_D_R_Z_R 0.1
`define AN4HSX4_C_F_Z_F 0.1
`define AN4HSX4_C_R_Z_R 0.1
`define AN4HSX4_B_F_Z_F 0.1
`define AN4HSX4_B_R_Z_R 0.1
`define AN4HSX4_A_F_Z_F 0.1
`define AN4HSX4_A_R_Z_R 0.1

module AN4HSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AN4HSX4_D_R_Z_R,`AN4HSX4_D_F_Z_F);
      (C +=> Z) = (`AN4HSX4_C_R_Z_R,`AN4HSX4_C_F_Z_F);
      (B +=> Z) = (`AN4HSX4_B_R_Z_R,`AN4HSX4_B_F_Z_F);
      (A +=> Z) = (`AN4HSX4_A_R_Z_R,`AN4HSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AN4HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:54 and Version :1.1 //

//  START
// CELL AN4HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN4HSX8_D_F_Z_F 0.1
`define AN4HSX8_D_R_Z_R 0.1
`define AN4HSX8_C_F_Z_F 0.1
`define AN4HSX8_C_R_Z_R 0.1
`define AN4HSX8_B_F_Z_F 0.1
`define AN4HSX8_B_R_Z_R 0.1
`define AN4HSX8_A_F_Z_F 0.1
`define AN4HSX8_A_R_Z_R 0.1

module AN4HSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AN4HSX8_D_R_Z_R,`AN4HSX8_D_F_Z_F);
      (C +=> Z) = (`AN4HSX8_C_R_Z_R,`AN4HSX8_C_F_Z_F);
      (B +=> Z) = (`AN4HSX8_B_R_Z_R,`AN4HSX8_B_F_Z_F);
      (A +=> Z) = (`AN4HSX8_A_R_Z_R,`AN4HSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AN4HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:02:54 and Version :1.1 //

//  START
// CELL AN5HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN5HS_E_F_Z_F 0.1
`define AN5HS_E_R_Z_R 0.1
`define AN5HS_D_F_Z_F 0.1
`define AN5HS_D_R_Z_R 0.1
`define AN5HS_C_F_Z_F 0.1
`define AN5HS_C_R_Z_R 0.1
`define AN5HS_B_F_Z_F 0.1
`define AN5HS_B_R_Z_R 0.1
`define AN5HS_A_F_Z_F 0.1
`define AN5HS_A_R_Z_R 0.1

module AN5HS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (Z, A, B, C, D, E);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AN5HS_E_R_Z_R,`AN5HS_E_F_Z_F);
      (D +=> Z) = (`AN5HS_D_R_Z_R,`AN5HS_D_F_Z_F);
      (C +=> Z) = (`AN5HS_C_R_Z_R,`AN5HS_C_F_Z_F);
      (B +=> Z) = (`AN5HS_B_R_Z_R,`AN5HS_B_F_Z_F);
      (A +=> Z) = (`AN5HS_A_R_Z_R,`AN5HS_A_F_Z_F);

   endspecify
`endif


endmodule // AN5HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:01 and Version :1.1 //
 
//  START 
// CELL AN5HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN5HSP_E_F_Z_F 0.1
`define AN5HSP_E_R_Z_R 0.1
`define AN5HSP_D_F_Z_F 0.1
`define AN5HSP_D_R_Z_R 0.1
`define AN5HSP_C_F_Z_F 0.1
`define AN5HSP_C_R_Z_R 0.1
`define AN5HSP_B_F_Z_F 0.1
`define AN5HSP_B_R_Z_R 0.1
`define AN5HSP_A_F_Z_F 0.1
`define AN5HSP_A_R_Z_R 0.1

module AN5HSP (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (Z, A, B, C, D, E);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AN5HSP_E_R_Z_R,`AN5HSP_E_F_Z_F);
      (D +=> Z) = (`AN5HSP_D_R_Z_R,`AN5HSP_D_F_Z_F);
      (C +=> Z) = (`AN5HSP_C_R_Z_R,`AN5HSP_C_F_Z_F);
      (B +=> Z) = (`AN5HSP_B_R_Z_R,`AN5HSP_B_F_Z_F);
      (A +=> Z) = (`AN5HSP_A_R_Z_R,`AN5HSP_A_F_Z_F);

   endspecify
`endif


endmodule // AN5HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:01 and Version :1.1 //
 
//  START 
// CELL AN5HSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN5HSX3_E_F_Z_F 0.1
`define AN5HSX3_E_R_Z_R 0.1
`define AN5HSX3_D_F_Z_F 0.1
`define AN5HSX3_D_R_Z_R 0.1
`define AN5HSX3_C_F_Z_F 0.1
`define AN5HSX3_C_R_Z_R 0.1
`define AN5HSX3_B_F_Z_F 0.1
`define AN5HSX3_B_R_Z_R 0.1
`define AN5HSX3_A_F_Z_F 0.1
`define AN5HSX3_A_R_Z_R 0.1

module AN5HSX3 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (Z, A, B, C, D, E);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AN5HSX3_E_R_Z_R,`AN5HSX3_E_F_Z_F);
      (D +=> Z) = (`AN5HSX3_D_R_Z_R,`AN5HSX3_D_F_Z_F);
      (C +=> Z) = (`AN5HSX3_C_R_Z_R,`AN5HSX3_C_F_Z_F);
      (B +=> Z) = (`AN5HSX3_B_R_Z_R,`AN5HSX3_B_F_Z_F);
      (A +=> Z) = (`AN5HSX3_A_R_Z_R,`AN5HSX3_A_F_Z_F);

   endspecify
`endif


endmodule // AN5HSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:01 and Version :1.1 //
 
//  START 
// CELL AN5HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN5HSX4_E_F_Z_F 0.1
`define AN5HSX4_E_R_Z_R 0.1
`define AN5HSX4_D_F_Z_F 0.1
`define AN5HSX4_D_R_Z_R 0.1
`define AN5HSX4_C_F_Z_F 0.1
`define AN5HSX4_C_R_Z_R 0.1
`define AN5HSX4_B_F_Z_F 0.1
`define AN5HSX4_B_R_Z_R 0.1
`define AN5HSX4_A_F_Z_F 0.1
`define AN5HSX4_A_R_Z_R 0.1

module AN5HSX4 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (Z, A, B, C, D, E);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AN5HSX4_E_R_Z_R,`AN5HSX4_E_F_Z_F);
      (D +=> Z) = (`AN5HSX4_D_R_Z_R,`AN5HSX4_D_F_Z_F);
      (C +=> Z) = (`AN5HSX4_C_R_Z_R,`AN5HSX4_C_F_Z_F);
      (B +=> Z) = (`AN5HSX4_B_R_Z_R,`AN5HSX4_B_F_Z_F);
      (A +=> Z) = (`AN5HSX4_A_R_Z_R,`AN5HSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AN5HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:01 and Version :1.1 //
 
//  START 
// CELL AN6HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN6HS_F_F_Z_F 0.1
`define AN6HS_F_R_Z_R 0.1
`define AN6HS_E_F_Z_F 0.1
`define AN6HS_E_R_Z_R 0.1
`define AN6HS_D_F_Z_F 0.1
`define AN6HS_D_R_Z_R 0.1
`define AN6HS_C_F_Z_F 0.1
`define AN6HS_C_R_Z_R 0.1
`define AN6HS_B_F_Z_F 0.1
`define AN6HS_B_R_Z_R 0.1
`define AN6HS_A_F_Z_F 0.1
`define AN6HS_A_R_Z_R 0.1

module AN6HS (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   and  u0 (Z, A, B, C, D, E, F);


`ifdef functional
`else
   specify

      (F +=> Z) = (`AN6HS_F_R_Z_R,`AN6HS_F_F_Z_F);
      (E +=> Z) = (`AN6HS_E_R_Z_R,`AN6HS_E_F_Z_F);
      (D +=> Z) = (`AN6HS_D_R_Z_R,`AN6HS_D_F_Z_F);
      (C +=> Z) = (`AN6HS_C_R_Z_R,`AN6HS_C_F_Z_F);
      (B +=> Z) = (`AN6HS_B_R_Z_R,`AN6HS_B_F_Z_F);
      (A +=> Z) = (`AN6HS_A_R_Z_R,`AN6HS_A_F_Z_F);

   endspecify
`endif


endmodule // AN6HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:04 and Version :1.1 //
 
//  START 
// CELL AN6HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN6HSP_F_F_Z_F 0.1
`define AN6HSP_F_R_Z_R 0.1
`define AN6HSP_E_F_Z_F 0.1
`define AN6HSP_E_R_Z_R 0.1
`define AN6HSP_D_F_Z_F 0.1
`define AN6HSP_D_R_Z_R 0.1
`define AN6HSP_C_F_Z_F 0.1
`define AN6HSP_C_R_Z_R 0.1
`define AN6HSP_B_F_Z_F 0.1
`define AN6HSP_B_R_Z_R 0.1
`define AN6HSP_A_F_Z_F 0.1
`define AN6HSP_A_R_Z_R 0.1

module AN6HSP (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   and  u0 (Z, A, B, C, D, E, F);


`ifdef functional
`else
   specify

      (F +=> Z) = (`AN6HSP_F_R_Z_R,`AN6HSP_F_F_Z_F);
      (E +=> Z) = (`AN6HSP_E_R_Z_R,`AN6HSP_E_F_Z_F);
      (D +=> Z) = (`AN6HSP_D_R_Z_R,`AN6HSP_D_F_Z_F);
      (C +=> Z) = (`AN6HSP_C_R_Z_R,`AN6HSP_C_F_Z_F);
      (B +=> Z) = (`AN6HSP_B_R_Z_R,`AN6HSP_B_F_Z_F);
      (A +=> Z) = (`AN6HSP_A_R_Z_R,`AN6HSP_A_F_Z_F);

   endspecify
`endif


endmodule // AN6HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:04 and Version :1.1 //
 
//  START 
// CELL AN6HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN6HSX4_F_F_Z_F 0.1
`define AN6HSX4_F_R_Z_R 0.1
`define AN6HSX4_E_F_Z_F 0.1
`define AN6HSX4_E_R_Z_R 0.1
`define AN6HSX4_D_F_Z_F 0.1
`define AN6HSX4_D_R_Z_R 0.1
`define AN6HSX4_C_F_Z_F 0.1
`define AN6HSX4_C_R_Z_R 0.1
`define AN6HSX4_B_F_Z_F 0.1
`define AN6HSX4_B_R_Z_R 0.1
`define AN6HSX4_A_F_Z_F 0.1
`define AN6HSX4_A_R_Z_R 0.1

module AN6HSX4 (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   and  u0 (Z, A, B, C, D, E, F);


`ifdef functional
`else
   specify

      (F +=> Z) = (`AN6HSX4_F_R_Z_R,`AN6HSX4_F_F_Z_F);
      (E +=> Z) = (`AN6HSX4_E_R_Z_R,`AN6HSX4_E_F_Z_F);
      (D +=> Z) = (`AN6HSX4_D_R_Z_R,`AN6HSX4_D_F_Z_F);
      (C +=> Z) = (`AN6HSX4_C_R_Z_R,`AN6HSX4_C_F_Z_F);
      (B +=> Z) = (`AN6HSX4_B_R_Z_R,`AN6HSX4_B_F_Z_F);
      (A +=> Z) = (`AN6HSX4_A_R_Z_R,`AN6HSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AN6HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:04 and Version :1.1 //
 
//  START 
// CELL AN7HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN7HS_G_F_Z_F 0.1
`define AN7HS_G_R_Z_R 0.1
`define AN7HS_F_F_Z_F 0.1
`define AN7HS_F_R_Z_R 0.1
`define AN7HS_E_F_Z_F 0.1
`define AN7HS_E_R_Z_R 0.1
`define AN7HS_D_F_Z_F 0.1
`define AN7HS_D_R_Z_R 0.1
`define AN7HS_C_F_Z_F 0.1
`define AN7HS_C_R_Z_R 0.1
`define AN7HS_B_F_Z_F 0.1
`define AN7HS_B_R_Z_R 0.1
`define AN7HS_A_F_Z_F 0.1
`define AN7HS_A_R_Z_R 0.1

module AN7HS (Z, A, B, C, D, E, F, G);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;
   input G;


   and  u0 (Z, A, B, C, D, E, F, G);


`ifdef functional
`else
   specify

      (G +=> Z) = (`AN7HS_G_R_Z_R,`AN7HS_G_F_Z_F);
      (F +=> Z) = (`AN7HS_F_R_Z_R,`AN7HS_F_F_Z_F);
      (E +=> Z) = (`AN7HS_E_R_Z_R,`AN7HS_E_F_Z_F);
      (D +=> Z) = (`AN7HS_D_R_Z_R,`AN7HS_D_F_Z_F);
      (C +=> Z) = (`AN7HS_C_R_Z_R,`AN7HS_C_F_Z_F);
      (B +=> Z) = (`AN7HS_B_R_Z_R,`AN7HS_B_F_Z_F);
      (A +=> Z) = (`AN7HS_A_R_Z_R,`AN7HS_A_F_Z_F);

   endspecify
`endif


endmodule // AN7HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:06 and Version :1.1 //
 
//  START 
// CELL AN7HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN7HSX4_G_F_Z_F 0.1
`define AN7HSX4_G_R_Z_R 0.1
`define AN7HSX4_F_F_Z_F 0.1
`define AN7HSX4_F_R_Z_R 0.1
`define AN7HSX4_E_F_Z_F 0.1
`define AN7HSX4_E_R_Z_R 0.1
`define AN7HSX4_D_F_Z_F 0.1
`define AN7HSX4_D_R_Z_R 0.1
`define AN7HSX4_C_F_Z_F 0.1
`define AN7HSX4_C_R_Z_R 0.1
`define AN7HSX4_B_F_Z_F 0.1
`define AN7HSX4_B_R_Z_R 0.1
`define AN7HSX4_A_F_Z_F 0.1
`define AN7HSX4_A_R_Z_R 0.1

module AN7HSX4 (Z, A, B, C, D, E, F, G);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;
   input G;


   and  u0 (Z, A, B, C, D, E, F, G);


`ifdef functional
`else
   specify

      (G +=> Z) = (`AN7HSX4_G_R_Z_R,`AN7HSX4_G_F_Z_F);
      (F +=> Z) = (`AN7HSX4_F_R_Z_R,`AN7HSX4_F_F_Z_F);
      (E +=> Z) = (`AN7HSX4_E_R_Z_R,`AN7HSX4_E_F_Z_F);
      (D +=> Z) = (`AN7HSX4_D_R_Z_R,`AN7HSX4_D_F_Z_F);
      (C +=> Z) = (`AN7HSX4_C_R_Z_R,`AN7HSX4_C_F_Z_F);
      (B +=> Z) = (`AN7HSX4_B_R_Z_R,`AN7HSX4_B_F_Z_F);
      (A +=> Z) = (`AN7HSX4_A_R_Z_R,`AN7HSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AN7HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:06 and Version :1.1 //
 
//  START 
// CELL AN8HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AN8HS_H_F_Z_F 0.1
`define AN8HS_H_R_Z_R 0.1
`define AN8HS_G_F_Z_F 0.1
`define AN8HS_G_R_Z_R 0.1
`define AN8HS_F_F_Z_F 0.1
`define AN8HS_F_R_Z_R 0.1
`define AN8HS_E_F_Z_F 0.1
`define AN8HS_E_R_Z_R 0.1
`define AN8HS_D_F_Z_F 0.1
`define AN8HS_D_R_Z_R 0.1
`define AN8HS_C_F_Z_F 0.1
`define AN8HS_C_R_Z_R 0.1
`define AN8HS_B_F_Z_F 0.1
`define AN8HS_B_R_Z_R 0.1
`define AN8HS_A_F_Z_F 0.1
`define AN8HS_A_R_Z_R 0.1

module AN8HS (Z, A, B, C, D, E, F, G, H);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;
   input G;
   input H;


   and  u0 (Z, A, B, C, D, E, F, G, H);


`ifdef functional
`else
   specify

      (H +=> Z) = (`AN8HS_H_R_Z_R,`AN8HS_H_F_Z_F);
      (G +=> Z) = (`AN8HS_G_R_Z_R,`AN8HS_G_F_Z_F);
      (F +=> Z) = (`AN8HS_F_R_Z_R,`AN8HS_F_F_Z_F);
      (E +=> Z) = (`AN8HS_E_R_Z_R,`AN8HS_E_F_Z_F);
      (D +=> Z) = (`AN8HS_D_R_Z_R,`AN8HS_D_F_Z_F);
      (C +=> Z) = (`AN8HS_C_R_Z_R,`AN8HS_C_F_Z_F);
      (B +=> Z) = (`AN8HS_B_R_Z_R,`AN8HS_B_F_Z_F);
      (A +=> Z) = (`AN8HS_A_R_Z_R,`AN8HS_A_F_Z_F);

   endspecify
`endif


endmodule // AN8HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:13 and Version :1.1 //
 
//  START 
// CELL AO1HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1HSX05_D_F_Z_R 0.1
`define AO1HSX05_D_R_Z_F 0.1
`define AO1HSX05_C_F_Z_R 0.1
`define AO1HSX05_C_R_Z_F 0.1
`define AO1HSX05_B_F_Z_R 0.1
`define AO1HSX05_B_R_Z_F 0.1
`define AO1HSX05_A_F_Z_R 0.1
`define AO1HSX05_A_R_Z_F 0.1

module AO1HSX05 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAB_, C, D);
   and  u1 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO1HSX05_D_F_Z_R,`AO1HSX05_D_R_Z_F);
      (C -=> Z) = (`AO1HSX05_C_F_Z_R,`AO1HSX05_C_R_Z_F);
      (B -=> Z) = (`AO1HSX05_B_F_Z_R,`AO1HSX05_B_R_Z_F);
      (A -=> Z) = (`AO1HSX05_A_F_Z_R,`AO1HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // AO1HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:15 and Version :1.1 //
 
//  START 
// CELL AO1HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1HS_D_F_Z_R 0.1
`define AO1HS_D_R_Z_F 0.1
`define AO1HS_C_F_Z_R 0.1
`define AO1HS_C_R_Z_F 0.1
`define AO1HS_B_F_Z_R 0.1
`define AO1HS_B_R_Z_F 0.1
`define AO1HS_A_F_Z_R 0.1
`define AO1HS_A_R_Z_F 0.1

module AO1HS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAB_, C, D);
   and  u1 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO1HS_D_F_Z_R,`AO1HS_D_R_Z_F);
      (C -=> Z) = (`AO1HS_C_F_Z_R,`AO1HS_C_R_Z_F);
      (B -=> Z) = (`AO1HS_B_F_Z_R,`AO1HS_B_R_Z_F);
      (A -=> Z) = (`AO1HS_A_F_Z_R,`AO1HS_A_R_Z_F);

   endspecify
`endif


endmodule // AO1HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:15 and Version :1.1 //
 
//  START 
// CELL AO1HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1HSP_D_F_Z_R 0.1
`define AO1HSP_D_R_Z_F 0.1
`define AO1HSP_C_F_Z_R 0.1
`define AO1HSP_C_R_Z_F 0.1
`define AO1HSP_B_F_Z_R 0.1
`define AO1HSP_B_R_Z_F 0.1
`define AO1HSP_A_F_Z_R 0.1
`define AO1HSP_A_R_Z_F 0.1

module AO1HSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAB_, C, D);
   and  u1 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO1HSP_D_F_Z_R,`AO1HSP_D_R_Z_F);
      (C -=> Z) = (`AO1HSP_C_F_Z_R,`AO1HSP_C_R_Z_F);
      (B -=> Z) = (`AO1HSP_B_F_Z_R,`AO1HSP_B_R_Z_F);
      (A -=> Z) = (`AO1HSP_A_F_Z_R,`AO1HSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO1HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:15 and Version :1.1 //
 
//  START 
// CELL AO1HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1HSX4_D_F_Z_R 0.1
`define AO1HSX4_D_R_Z_F 0.1
`define AO1HSX4_C_F_Z_R 0.1
`define AO1HSX4_C_R_Z_F 0.1
`define AO1HSX4_B_F_Z_R 0.1
`define AO1HSX4_B_R_Z_F 0.1
`define AO1HSX4_A_F_Z_R 0.1
`define AO1HSX4_A_R_Z_F 0.1

module AO1HSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAB_, C, D);
   and  u1 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO1HSX4_D_F_Z_R,`AO1HSX4_D_R_Z_F);
      (C -=> Z) = (`AO1HSX4_C_F_Z_R,`AO1HSX4_C_R_Z_F);
      (B -=> Z) = (`AO1HSX4_B_F_Z_R,`AO1HSX4_B_R_Z_F);
      (A -=> Z) = (`AO1HSX4_A_F_Z_R,`AO1HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO1HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:15 and Version :1.1 //
 
//  START 
// CELL AO1HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1HSX8_D_F_Z_R 0.1
`define AO1HSX8_D_R_Z_F 0.1
`define AO1HSX8_C_F_Z_R 0.1
`define AO1HSX8_C_R_Z_F 0.1
`define AO1HSX8_B_F_Z_R 0.1
`define AO1HSX8_B_R_Z_F 0.1
`define AO1HSX8_A_F_Z_R 0.1
`define AO1HSX8_A_R_Z_F 0.1

module AO1HSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAB_, C, D);
   and  u1 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO1HSX8_D_F_Z_R,`AO1HSX8_D_R_Z_F);
      (C -=> Z) = (`AO1HSX8_C_F_Z_R,`AO1HSX8_C_R_Z_F);
      (B -=> Z) = (`AO1HSX8_B_F_Z_R,`AO1HSX8_B_R_Z_F);
      (A -=> Z) = (`AO1HSX8_A_F_Z_R,`AO1HSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AO1HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:15 and Version :1.1 //
 
//  START 
// CELL AO10HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO10HSX05_E_F_Z_R 0.1
`define AO10HSX05_E_R_Z_F 0.1
`define AO10HSX05_D_F_Z_R 0.1
`define AO10HSX05_D_R_Z_F 0.1
`define AO10HSX05_C_F_Z_R 0.1
`define AO10HSX05_C_R_Z_F 0.1
`define AO10HSX05_B_F_Z_R 0.1
`define AO10HSX05_B_R_Z_F 0.1
`define AO10HSX05_A_F_Z_R 0.1
`define AO10HSX05_A_R_Z_F 0.1

module AO10HSX05 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   nor  u0 (Z, AndAB_, AndCD_, E);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (E -=> Z) = (`AO10HSX05_E_F_Z_R,`AO10HSX05_E_R_Z_F);
      (D -=> Z) = (`AO10HSX05_D_F_Z_R,`AO10HSX05_D_R_Z_F);
      (C -=> Z) = (`AO10HSX05_C_F_Z_R,`AO10HSX05_C_R_Z_F);
      (B -=> Z) = (`AO10HSX05_B_F_Z_R,`AO10HSX05_B_R_Z_F);
      (A -=> Z) = (`AO10HSX05_A_F_Z_R,`AO10HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // AO10HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:31 and Version :1.1 //
 
//  START 
// CELL AO10HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO10HS_E_F_Z_R 0.1
`define AO10HS_E_R_Z_F 0.1
`define AO10HS_D_F_Z_R 0.1
`define AO10HS_D_R_Z_F 0.1
`define AO10HS_C_F_Z_R 0.1
`define AO10HS_C_R_Z_F 0.1
`define AO10HS_B_F_Z_R 0.1
`define AO10HS_B_R_Z_F 0.1
`define AO10HS_A_F_Z_R 0.1
`define AO10HS_A_R_Z_F 0.1

module AO10HS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   nor  u0 (Z, AndAB_, AndCD_, E);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (E -=> Z) = (`AO10HS_E_F_Z_R,`AO10HS_E_R_Z_F);
      (D -=> Z) = (`AO10HS_D_F_Z_R,`AO10HS_D_R_Z_F);
      (C -=> Z) = (`AO10HS_C_F_Z_R,`AO10HS_C_R_Z_F);
      (B -=> Z) = (`AO10HS_B_F_Z_R,`AO10HS_B_R_Z_F);
      (A -=> Z) = (`AO10HS_A_F_Z_R,`AO10HS_A_R_Z_F);

   endspecify
`endif


endmodule // AO10HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:31 and Version :1.1 //
 
//  START 
// CELL AO10HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO10HSP_E_F_Z_R 0.1
`define AO10HSP_E_R_Z_F 0.1
`define AO10HSP_D_F_Z_R 0.1
`define AO10HSP_D_R_Z_F 0.1
`define AO10HSP_C_F_Z_R 0.1
`define AO10HSP_C_R_Z_F 0.1
`define AO10HSP_B_F_Z_R 0.1
`define AO10HSP_B_R_Z_F 0.1
`define AO10HSP_A_F_Z_R 0.1
`define AO10HSP_A_R_Z_F 0.1

module AO10HSP (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   nor  u0 (Z, AndAB_, AndCD_, E);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (E -=> Z) = (`AO10HSP_E_F_Z_R,`AO10HSP_E_R_Z_F);
      (D -=> Z) = (`AO10HSP_D_F_Z_R,`AO10HSP_D_R_Z_F);
      (C -=> Z) = (`AO10HSP_C_F_Z_R,`AO10HSP_C_R_Z_F);
      (B -=> Z) = (`AO10HSP_B_F_Z_R,`AO10HSP_B_R_Z_F);
      (A -=> Z) = (`AO10HSP_A_F_Z_R,`AO10HSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO10HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:31 and Version :1.1 //
 
//  START 
// CELL AO10HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO10HSX4_E_F_Z_R 0.1
`define AO10HSX4_E_R_Z_F 0.1
`define AO10HSX4_D_F_Z_R 0.1
`define AO10HSX4_D_R_Z_F 0.1
`define AO10HSX4_C_F_Z_R 0.1
`define AO10HSX4_C_R_Z_F 0.1
`define AO10HSX4_B_F_Z_R 0.1
`define AO10HSX4_B_R_Z_F 0.1
`define AO10HSX4_A_F_Z_R 0.1
`define AO10HSX4_A_R_Z_F 0.1

module AO10HSX4 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   nor  u0 (Z, AndAB_, AndCD_, E);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (E -=> Z) = (`AO10HSX4_E_F_Z_R,`AO10HSX4_E_R_Z_F);
      (D -=> Z) = (`AO10HSX4_D_F_Z_R,`AO10HSX4_D_R_Z_F);
      (C -=> Z) = (`AO10HSX4_C_F_Z_R,`AO10HSX4_C_R_Z_F);
      (B -=> Z) = (`AO10HSX4_B_F_Z_R,`AO10HSX4_B_R_Z_F);
      (A -=> Z) = (`AO10HSX4_A_F_Z_R,`AO10HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO10HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:31 and Version :1.1 //
 
//  START 
// CELL AO10HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO10HSX8_E_F_Z_R 0.1
`define AO10HSX8_E_R_Z_F 0.1
`define AO10HSX8_D_F_Z_R 0.1
`define AO10HSX8_D_R_Z_F 0.1
`define AO10HSX8_C_F_Z_R 0.1
`define AO10HSX8_C_R_Z_F 0.1
`define AO10HSX8_B_F_Z_R 0.1
`define AO10HSX8_B_R_Z_F 0.1
`define AO10HSX8_A_F_Z_R 0.1
`define AO10HSX8_A_R_Z_F 0.1

module AO10HSX8 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   nor  u0 (Z, AndAB_, AndCD_, E);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (E -=> Z) = (`AO10HSX8_E_F_Z_R,`AO10HSX8_E_R_Z_F);
      (D -=> Z) = (`AO10HSX8_D_F_Z_R,`AO10HSX8_D_R_Z_F);
      (C -=> Z) = (`AO10HSX8_C_F_Z_R,`AO10HSX8_C_R_Z_F);
      (B -=> Z) = (`AO10HSX8_B_F_Z_R,`AO10HSX8_B_R_Z_F);
      (A -=> Z) = (`AO10HSX8_A_F_Z_R,`AO10HSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AO10HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:31 and Version :1.1 //
 
//  START 
// CELL AO10NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO10NHS_E_F_Z_F 0.1
`define AO10NHS_E_R_Z_R 0.1
`define AO10NHS_D_F_Z_F 0.1
`define AO10NHS_D_R_Z_R 0.1
`define AO10NHS_C_F_Z_F 0.1
`define AO10NHS_C_R_Z_R 0.1
`define AO10NHS_B_F_Z_F 0.1
`define AO10NHS_B_R_Z_R 0.1
`define AO10NHS_A_F_Z_F 0.1
`define AO10NHS_A_R_Z_R 0.1

module AO10NHS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndAB_, A, B);
   and  u1 (AndCD_, C, D);
   or  u2 (Z, AndAB_, AndCD_, E);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO10NHS_E_R_Z_R,`AO10NHS_E_F_Z_F);
      (D +=> Z) = (`AO10NHS_D_R_Z_R,`AO10NHS_D_F_Z_F);
      (C +=> Z) = (`AO10NHS_C_R_Z_R,`AO10NHS_C_F_Z_F);
      (B +=> Z) = (`AO10NHS_B_R_Z_R,`AO10NHS_B_F_Z_F);
      (A +=> Z) = (`AO10NHS_A_R_Z_R,`AO10NHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO10NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:31 and Version :1.1 //
 
//  START 
// CELL AO10NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO10NHSP_E_F_Z_F 0.1
`define AO10NHSP_E_R_Z_R 0.1
`define AO10NHSP_D_F_Z_F 0.1
`define AO10NHSP_D_R_Z_R 0.1
`define AO10NHSP_C_F_Z_F 0.1
`define AO10NHSP_C_R_Z_R 0.1
`define AO10NHSP_B_F_Z_F 0.1
`define AO10NHSP_B_R_Z_R 0.1
`define AO10NHSP_A_F_Z_F 0.1
`define AO10NHSP_A_R_Z_R 0.1

module AO10NHSP (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndAB_, A, B);
   and  u1 (AndCD_, C, D);
   or  u2 (Z, AndAB_, AndCD_, E);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO10NHSP_E_R_Z_R,`AO10NHSP_E_F_Z_F);
      (D +=> Z) = (`AO10NHSP_D_R_Z_R,`AO10NHSP_D_F_Z_F);
      (C +=> Z) = (`AO10NHSP_C_R_Z_R,`AO10NHSP_C_F_Z_F);
      (B +=> Z) = (`AO10NHSP_B_R_Z_R,`AO10NHSP_B_F_Z_F);
      (A +=> Z) = (`AO10NHSP_A_R_Z_R,`AO10NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO10NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:31 and Version :1.1 //
 
//  START 
// CELL AO10NHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO10NHSX4_E_F_Z_F 0.1
`define AO10NHSX4_E_R_Z_R 0.1
`define AO10NHSX4_D_F_Z_F 0.1
`define AO10NHSX4_D_R_Z_R 0.1
`define AO10NHSX4_C_F_Z_F 0.1
`define AO10NHSX4_C_R_Z_R 0.1
`define AO10NHSX4_B_F_Z_F 0.1
`define AO10NHSX4_B_R_Z_R 0.1
`define AO10NHSX4_A_F_Z_F 0.1
`define AO10NHSX4_A_R_Z_R 0.1

module AO10NHSX4 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndAB_, A, B);
   and  u1 (AndCD_, C, D);
   or  u2 (Z, AndAB_, AndCD_, E);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO10NHSX4_E_R_Z_R,`AO10NHSX4_E_F_Z_F);
      (D +=> Z) = (`AO10NHSX4_D_R_Z_R,`AO10NHSX4_D_F_Z_F);
      (C +=> Z) = (`AO10NHSX4_C_R_Z_R,`AO10NHSX4_C_F_Z_F);
      (B +=> Z) = (`AO10NHSX4_B_R_Z_R,`AO10NHSX4_B_F_Z_F);
      (A +=> Z) = (`AO10NHSX4_A_R_Z_R,`AO10NHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO10NHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:31 and Version :1.1 //
 
//  START 
// CELL AO10NHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO10NHSX8_E_F_Z_F 0.1
`define AO10NHSX8_E_R_Z_R 0.1
`define AO10NHSX8_D_F_Z_F 0.1
`define AO10NHSX8_D_R_Z_R 0.1
`define AO10NHSX8_C_F_Z_F 0.1
`define AO10NHSX8_C_R_Z_R 0.1
`define AO10NHSX8_B_F_Z_F 0.1
`define AO10NHSX8_B_R_Z_R 0.1
`define AO10NHSX8_A_F_Z_F 0.1
`define AO10NHSX8_A_R_Z_R 0.1

module AO10NHSX8 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndAB_, A, B);
   and  u1 (AndCD_, C, D);
   or  u2 (Z, AndAB_, AndCD_, E);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO10NHSX8_E_R_Z_R,`AO10NHSX8_E_F_Z_F);
      (D +=> Z) = (`AO10NHSX8_D_R_Z_R,`AO10NHSX8_D_F_Z_F);
      (C +=> Z) = (`AO10NHSX8_C_R_Z_R,`AO10NHSX8_C_F_Z_F);
      (B +=> Z) = (`AO10NHSX8_B_R_Z_R,`AO10NHSX8_B_F_Z_F);
      (A +=> Z) = (`AO10NHSX8_A_R_Z_R,`AO10NHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO10NHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:31 and Version :1.1 //
 
//  START 
// CELL F_AO10NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO10NHS_E_F_Z_F 0.1
`define F_AO10NHS_E_R_Z_R 0.1
`define F_AO10NHS_D_F_Z_F 0.1
`define F_AO10NHS_D_R_Z_R 0.1
`define F_AO10NHS_C_F_Z_F 0.1
`define F_AO10NHS_C_R_Z_R 0.1
`define F_AO10NHS_B_F_Z_F 0.1
`define F_AO10NHS_B_R_Z_R 0.1
`define F_AO10NHS_A_F_Z_F 0.1
`define F_AO10NHS_A_R_Z_R 0.1

module F_AO10NHS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndAB_, A, B);
   and  u1 (AndCD_, C, D);
   or  u2 (Z, AndAB_, AndCD_, E);


`ifdef functional
`else
   specify

      (E +=> Z) = (`F_AO10NHS_E_R_Z_R,`F_AO10NHS_E_F_Z_F);
      (D +=> Z) = (`F_AO10NHS_D_R_Z_R,`F_AO10NHS_D_F_Z_F);
      (C +=> Z) = (`F_AO10NHS_C_R_Z_R,`F_AO10NHS_C_F_Z_F);
      (B +=> Z) = (`F_AO10NHS_B_R_Z_R,`F_AO10NHS_B_F_Z_F);
      (A +=> Z) = (`F_AO10NHS_A_R_Z_R,`F_AO10NHS_A_F_Z_F);

   endspecify
`endif


endmodule // F_AO10NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:31 and Version :1.1 //
 
//  START 
// CELL F_AO10NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO10NHSP_E_F_Z_F 0.1
`define F_AO10NHSP_E_R_Z_R 0.1
`define F_AO10NHSP_D_F_Z_F 0.1
`define F_AO10NHSP_D_R_Z_R 0.1
`define F_AO10NHSP_C_F_Z_F 0.1
`define F_AO10NHSP_C_R_Z_R 0.1
`define F_AO10NHSP_B_F_Z_F 0.1
`define F_AO10NHSP_B_R_Z_R 0.1
`define F_AO10NHSP_A_F_Z_F 0.1
`define F_AO10NHSP_A_R_Z_R 0.1

module F_AO10NHSP (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndAB_, A, B);
   and  u1 (AndCD_, C, D);
   or  u2 (Z, AndAB_, AndCD_, E);


`ifdef functional
`else
   specify

      (E +=> Z) = (`F_AO10NHSP_E_R_Z_R,`F_AO10NHSP_E_F_Z_F);
      (D +=> Z) = (`F_AO10NHSP_D_R_Z_R,`F_AO10NHSP_D_F_Z_F);
      (C +=> Z) = (`F_AO10NHSP_C_R_Z_R,`F_AO10NHSP_C_F_Z_F);
      (B +=> Z) = (`F_AO10NHSP_B_R_Z_R,`F_AO10NHSP_B_F_Z_F);
      (A +=> Z) = (`F_AO10NHSP_A_R_Z_R,`F_AO10NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // F_AO10NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:31 and Version :1.1 //
 
//  START 
// CELL AO11HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO11HSX05_F_F_Z_R 0.1
`define AO11HSX05_F_R_Z_F 0.1
`define AO11HSX05_E_F_Z_R 0.1
`define AO11HSX05_E_R_Z_F 0.1
`define AO11HSX05_D_F_Z_R 0.1
`define AO11HSX05_D_R_Z_F 0.1
`define AO11HSX05_C_F_Z_R 0.1
`define AO11HSX05_C_R_Z_F 0.1
`define AO11HSX05_B_F_Z_R 0.1
`define AO11HSX05_B_R_Z_F 0.1
`define AO11HSX05_A_F_Z_R 0.1
`define AO11HSX05_A_R_Z_F 0.1

module AO11HSX05 (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   nor  u0 (Z, AndAB_, AndCD_, AndEF_);
   and  u1 (AndEF_, E, F);
   and  u2 (AndCD_, C, D);
   and  u3 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (F -=> Z) = (`AO11HSX05_F_F_Z_R,`AO11HSX05_F_R_Z_F);
      (E -=> Z) = (`AO11HSX05_E_F_Z_R,`AO11HSX05_E_R_Z_F);
      (D -=> Z) = (`AO11HSX05_D_F_Z_R,`AO11HSX05_D_R_Z_F);
      (C -=> Z) = (`AO11HSX05_C_F_Z_R,`AO11HSX05_C_R_Z_F);
      (B -=> Z) = (`AO11HSX05_B_F_Z_R,`AO11HSX05_B_R_Z_F);
      (A -=> Z) = (`AO11HSX05_A_F_Z_R,`AO11HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // AO11HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:43 and Version :1.1 //
 
//  START 
// CELL AO11HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO11HS_F_F_Z_R 0.1
`define AO11HS_F_R_Z_F 0.1
`define AO11HS_E_F_Z_R 0.1
`define AO11HS_E_R_Z_F 0.1
`define AO11HS_D_F_Z_R 0.1
`define AO11HS_D_R_Z_F 0.1
`define AO11HS_C_F_Z_R 0.1
`define AO11HS_C_R_Z_F 0.1
`define AO11HS_B_F_Z_R 0.1
`define AO11HS_B_R_Z_F 0.1
`define AO11HS_A_F_Z_R 0.1
`define AO11HS_A_R_Z_F 0.1

module AO11HS (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   nor  u0 (Z, AndAB_, AndCD_, AndEF_);
   and  u1 (AndEF_, E, F);
   and  u2 (AndCD_, C, D);
   and  u3 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (F -=> Z) = (`AO11HS_F_F_Z_R,`AO11HS_F_R_Z_F);
      (E -=> Z) = (`AO11HS_E_F_Z_R,`AO11HS_E_R_Z_F);
      (D -=> Z) = (`AO11HS_D_F_Z_R,`AO11HS_D_R_Z_F);
      (C -=> Z) = (`AO11HS_C_F_Z_R,`AO11HS_C_R_Z_F);
      (B -=> Z) = (`AO11HS_B_F_Z_R,`AO11HS_B_R_Z_F);
      (A -=> Z) = (`AO11HS_A_F_Z_R,`AO11HS_A_R_Z_F);

   endspecify
`endif


endmodule // AO11HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:43 and Version :1.1 //
 
//  START 
// CELL AO11HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO11HSP_F_F_Z_R 0.1
`define AO11HSP_F_R_Z_F 0.1
`define AO11HSP_E_F_Z_R 0.1
`define AO11HSP_E_R_Z_F 0.1
`define AO11HSP_D_F_Z_R 0.1
`define AO11HSP_D_R_Z_F 0.1
`define AO11HSP_C_F_Z_R 0.1
`define AO11HSP_C_R_Z_F 0.1
`define AO11HSP_B_F_Z_R 0.1
`define AO11HSP_B_R_Z_F 0.1
`define AO11HSP_A_F_Z_R 0.1
`define AO11HSP_A_R_Z_F 0.1

module AO11HSP (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   nor  u0 (Z, AndAB_, AndCD_, AndEF_);
   and  u1 (AndEF_, E, F);
   and  u2 (AndCD_, C, D);
   and  u3 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (F -=> Z) = (`AO11HSP_F_F_Z_R,`AO11HSP_F_R_Z_F);
      (E -=> Z) = (`AO11HSP_E_F_Z_R,`AO11HSP_E_R_Z_F);
      (D -=> Z) = (`AO11HSP_D_F_Z_R,`AO11HSP_D_R_Z_F);
      (C -=> Z) = (`AO11HSP_C_F_Z_R,`AO11HSP_C_R_Z_F);
      (B -=> Z) = (`AO11HSP_B_F_Z_R,`AO11HSP_B_R_Z_F);
      (A -=> Z) = (`AO11HSP_A_F_Z_R,`AO11HSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO11HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:43 and Version :1.1 //
 
//  START 
// CELL AO11HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO11HSX4_F_F_Z_R 0.1
`define AO11HSX4_F_R_Z_F 0.1
`define AO11HSX4_E_F_Z_R 0.1
`define AO11HSX4_E_R_Z_F 0.1
`define AO11HSX4_D_F_Z_R 0.1
`define AO11HSX4_D_R_Z_F 0.1
`define AO11HSX4_C_F_Z_R 0.1
`define AO11HSX4_C_R_Z_F 0.1
`define AO11HSX4_B_F_Z_R 0.1
`define AO11HSX4_B_R_Z_F 0.1
`define AO11HSX4_A_F_Z_R 0.1
`define AO11HSX4_A_R_Z_F 0.1

module AO11HSX4 (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   nor  u0 (Z, AndAB_, AndCD_, AndEF_);
   and  u1 (AndEF_, E, F);
   and  u2 (AndCD_, C, D);
   and  u3 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (F -=> Z) = (`AO11HSX4_F_F_Z_R,`AO11HSX4_F_R_Z_F);
      (E -=> Z) = (`AO11HSX4_E_F_Z_R,`AO11HSX4_E_R_Z_F);
      (D -=> Z) = (`AO11HSX4_D_F_Z_R,`AO11HSX4_D_R_Z_F);
      (C -=> Z) = (`AO11HSX4_C_F_Z_R,`AO11HSX4_C_R_Z_F);
      (B -=> Z) = (`AO11HSX4_B_F_Z_R,`AO11HSX4_B_R_Z_F);
      (A -=> Z) = (`AO11HSX4_A_F_Z_R,`AO11HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO11HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:43 and Version :1.1 //
 
//  START 
// CELL AO11HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO11HSX8_F_F_Z_R 0.1
`define AO11HSX8_F_R_Z_F 0.1
`define AO11HSX8_E_F_Z_R 0.1
`define AO11HSX8_E_R_Z_F 0.1
`define AO11HSX8_D_F_Z_R 0.1
`define AO11HSX8_D_R_Z_F 0.1
`define AO11HSX8_C_F_Z_R 0.1
`define AO11HSX8_C_R_Z_F 0.1
`define AO11HSX8_B_F_Z_R 0.1
`define AO11HSX8_B_R_Z_F 0.1
`define AO11HSX8_A_F_Z_R 0.1
`define AO11HSX8_A_R_Z_F 0.1

module AO11HSX8 (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   nor  u0 (Z, AndAB_, AndCD_, AndEF_);
   and  u1 (AndEF_, E, F);
   and  u2 (AndCD_, C, D);
   and  u3 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (F -=> Z) = (`AO11HSX8_F_F_Z_R,`AO11HSX8_F_R_Z_F);
      (E -=> Z) = (`AO11HSX8_E_F_Z_R,`AO11HSX8_E_R_Z_F);
      (D -=> Z) = (`AO11HSX8_D_F_Z_R,`AO11HSX8_D_R_Z_F);
      (C -=> Z) = (`AO11HSX8_C_F_Z_R,`AO11HSX8_C_R_Z_F);
      (B -=> Z) = (`AO11HSX8_B_F_Z_R,`AO11HSX8_B_R_Z_F);
      (A -=> Z) = (`AO11HSX8_A_F_Z_R,`AO11HSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AO11HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:43 and Version :1.1 //
 
//  START 
// CELL AO11NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO11NHS_F_F_Z_F 0.1
`define AO11NHS_F_R_Z_R 0.1
`define AO11NHS_E_F_Z_F 0.1
`define AO11NHS_E_R_Z_R 0.1
`define AO11NHS_D_F_Z_F 0.1
`define AO11NHS_D_R_Z_R 0.1
`define AO11NHS_C_F_Z_F 0.1
`define AO11NHS_C_R_Z_R 0.1
`define AO11NHS_B_F_Z_F 0.1
`define AO11NHS_B_R_Z_R 0.1
`define AO11NHS_A_F_Z_F 0.1
`define AO11NHS_A_R_Z_R 0.1

module AO11NHS (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   and  u0 (AndAB_, A, B);
   and  u1 (AndCD_, C, D);
   and  u2 (AndEF_, E, F);
   or  u3 (Z, AndAB_, AndCD_, AndEF_);


`ifdef functional
`else
   specify

      (F +=> Z) = (`AO11NHS_F_R_Z_R,`AO11NHS_F_F_Z_F);
      (E +=> Z) = (`AO11NHS_E_R_Z_R,`AO11NHS_E_F_Z_F);
      (D +=> Z) = (`AO11NHS_D_R_Z_R,`AO11NHS_D_F_Z_F);
      (C +=> Z) = (`AO11NHS_C_R_Z_R,`AO11NHS_C_F_Z_F);
      (B +=> Z) = (`AO11NHS_B_R_Z_R,`AO11NHS_B_F_Z_F);
      (A +=> Z) = (`AO11NHS_A_R_Z_R,`AO11NHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO11NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:43 and Version :1.1 //
 
//  START 
// CELL AO11NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO11NHSP_F_F_Z_F 0.1
`define AO11NHSP_F_R_Z_R 0.1
`define AO11NHSP_E_F_Z_F 0.1
`define AO11NHSP_E_R_Z_R 0.1
`define AO11NHSP_D_F_Z_F 0.1
`define AO11NHSP_D_R_Z_R 0.1
`define AO11NHSP_C_F_Z_F 0.1
`define AO11NHSP_C_R_Z_R 0.1
`define AO11NHSP_B_F_Z_F 0.1
`define AO11NHSP_B_R_Z_R 0.1
`define AO11NHSP_A_F_Z_F 0.1
`define AO11NHSP_A_R_Z_R 0.1

module AO11NHSP (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   and  u0 (AndAB_, A, B);
   and  u1 (AndCD_, C, D);
   and  u2 (AndEF_, E, F);
   or  u3 (Z, AndAB_, AndCD_, AndEF_);


`ifdef functional
`else
   specify

      (F +=> Z) = (`AO11NHSP_F_R_Z_R,`AO11NHSP_F_F_Z_F);
      (E +=> Z) = (`AO11NHSP_E_R_Z_R,`AO11NHSP_E_F_Z_F);
      (D +=> Z) = (`AO11NHSP_D_R_Z_R,`AO11NHSP_D_F_Z_F);
      (C +=> Z) = (`AO11NHSP_C_R_Z_R,`AO11NHSP_C_F_Z_F);
      (B +=> Z) = (`AO11NHSP_B_R_Z_R,`AO11NHSP_B_F_Z_F);
      (A +=> Z) = (`AO11NHSP_A_R_Z_R,`AO11NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO11NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:43 and Version :1.1 //
 
//  START 
// CELL AO11NHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO11NHSX4_F_F_Z_F 0.1
`define AO11NHSX4_F_R_Z_R 0.1
`define AO11NHSX4_E_F_Z_F 0.1
`define AO11NHSX4_E_R_Z_R 0.1
`define AO11NHSX4_D_F_Z_F 0.1
`define AO11NHSX4_D_R_Z_R 0.1
`define AO11NHSX4_C_F_Z_F 0.1
`define AO11NHSX4_C_R_Z_R 0.1
`define AO11NHSX4_B_F_Z_F 0.1
`define AO11NHSX4_B_R_Z_R 0.1
`define AO11NHSX4_A_F_Z_F 0.1
`define AO11NHSX4_A_R_Z_R 0.1

module AO11NHSX4 (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   and  u0 (AndAB_, A, B);
   and  u1 (AndCD_, C, D);
   and  u2 (AndEF_, E, F);
   or  u3 (Z, AndAB_, AndCD_, AndEF_);


`ifdef functional
`else
   specify

      (F +=> Z) = (`AO11NHSX4_F_R_Z_R,`AO11NHSX4_F_F_Z_F);
      (E +=> Z) = (`AO11NHSX4_E_R_Z_R,`AO11NHSX4_E_F_Z_F);
      (D +=> Z) = (`AO11NHSX4_D_R_Z_R,`AO11NHSX4_D_F_Z_F);
      (C +=> Z) = (`AO11NHSX4_C_R_Z_R,`AO11NHSX4_C_F_Z_F);
      (B +=> Z) = (`AO11NHSX4_B_R_Z_R,`AO11NHSX4_B_F_Z_F);
      (A +=> Z) = (`AO11NHSX4_A_R_Z_R,`AO11NHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO11NHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:43 and Version :1.1 //
 
//  START 
// CELL AO11NHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO11NHSX8_F_F_Z_F 0.1
`define AO11NHSX8_F_R_Z_R 0.1
`define AO11NHSX8_E_F_Z_F 0.1
`define AO11NHSX8_E_R_Z_R 0.1
`define AO11NHSX8_D_F_Z_F 0.1
`define AO11NHSX8_D_R_Z_R 0.1
`define AO11NHSX8_C_F_Z_F 0.1
`define AO11NHSX8_C_R_Z_R 0.1
`define AO11NHSX8_B_F_Z_F 0.1
`define AO11NHSX8_B_R_Z_R 0.1
`define AO11NHSX8_A_F_Z_F 0.1
`define AO11NHSX8_A_R_Z_R 0.1

module AO11NHSX8 (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   and  u0 (AndAB_, A, B);
   and  u1 (AndCD_, C, D);
   and  u2 (AndEF_, E, F);
   or  u3 (Z, AndAB_, AndCD_, AndEF_);


`ifdef functional
`else
   specify

      (F +=> Z) = (`AO11NHSX8_F_R_Z_R,`AO11NHSX8_F_F_Z_F);
      (E +=> Z) = (`AO11NHSX8_E_R_Z_R,`AO11NHSX8_E_F_Z_F);
      (D +=> Z) = (`AO11NHSX8_D_R_Z_R,`AO11NHSX8_D_F_Z_F);
      (C +=> Z) = (`AO11NHSX8_C_R_Z_R,`AO11NHSX8_C_F_Z_F);
      (B +=> Z) = (`AO11NHSX8_B_R_Z_R,`AO11NHSX8_B_F_Z_F);
      (A +=> Z) = (`AO11NHSX8_A_R_Z_R,`AO11NHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO11NHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:43 and Version :1.1 //
 
//  START 
// CELL F_AO11NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO11NHSP_F_F_Z_F 0.1
`define F_AO11NHSP_F_R_Z_R 0.1
`define F_AO11NHSP_E_F_Z_F 0.1
`define F_AO11NHSP_E_R_Z_R 0.1
`define F_AO11NHSP_D_F_Z_F 0.1
`define F_AO11NHSP_D_R_Z_R 0.1
`define F_AO11NHSP_C_F_Z_F 0.1
`define F_AO11NHSP_C_R_Z_R 0.1
`define F_AO11NHSP_B_F_Z_F 0.1
`define F_AO11NHSP_B_R_Z_R 0.1
`define F_AO11NHSP_A_F_Z_F 0.1
`define F_AO11NHSP_A_R_Z_R 0.1

module F_AO11NHSP (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   and  u0 (AndAB_, A, B);
   and  u1 (AndCD_, C, D);
   and  u2 (AndEF_, E, F);
   or  u3 (Z, AndAB_, AndCD_, AndEF_);


`ifdef functional
`else
   specify

      (F +=> Z) = (`F_AO11NHSP_F_R_Z_R,`F_AO11NHSP_F_F_Z_F);
      (E +=> Z) = (`F_AO11NHSP_E_R_Z_R,`F_AO11NHSP_E_F_Z_F);
      (D +=> Z) = (`F_AO11NHSP_D_R_Z_R,`F_AO11NHSP_D_F_Z_F);
      (C +=> Z) = (`F_AO11NHSP_C_R_Z_R,`F_AO11NHSP_C_F_Z_F);
      (B +=> Z) = (`F_AO11NHSP_B_R_Z_R,`F_AO11NHSP_B_F_Z_F);
      (A +=> Z) = (`F_AO11NHSP_A_R_Z_R,`F_AO11NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // F_AO11NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:43 and Version :1.1 //
 
//  START 
// CELL AO12HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO12HS_H_F_Z_R 0.1
`define AO12HS_H_R_Z_F 0.1
`define AO12HS_G_F_Z_R 0.1
`define AO12HS_G_R_Z_F 0.1
`define AO12HS_F_F_Z_R 0.1
`define AO12HS_F_R_Z_F 0.1
`define AO12HS_E_F_Z_R 0.1
`define AO12HS_E_R_Z_F 0.1
`define AO12HS_D_F_Z_R 0.1
`define AO12HS_D_R_Z_F 0.1
`define AO12HS_C_F_Z_R 0.1
`define AO12HS_C_R_Z_F 0.1
`define AO12HS_B_F_Z_R 0.1
`define AO12HS_B_R_Z_F 0.1
`define AO12HS_A_F_Z_R 0.1
`define AO12HS_A_R_Z_F 0.1

module AO12HS (Z, A, B, C, D, E, F, G, H);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;
   input G;
   input H;


   or  u0 (OrAB_, A, B);
   or  u1 (OrCD_, C, D);
   or  u2 (OrEF_, E, F);
   or  u3 (OrGH_, G, H);
   nand  u4 (Z, OrAB_, OrCD_, OrEF_, OrGH_);


`ifdef functional
`else
   specify

      (H -=> Z) = (`AO12HS_H_F_Z_R,`AO12HS_H_R_Z_F);
      (G -=> Z) = (`AO12HS_G_F_Z_R,`AO12HS_G_R_Z_F);
      (F -=> Z) = (`AO12HS_F_F_Z_R,`AO12HS_F_R_Z_F);
      (E -=> Z) = (`AO12HS_E_F_Z_R,`AO12HS_E_R_Z_F);
      (D -=> Z) = (`AO12HS_D_F_Z_R,`AO12HS_D_R_Z_F);
      (C -=> Z) = (`AO12HS_C_F_Z_R,`AO12HS_C_R_Z_F);
      (B -=> Z) = (`AO12HS_B_F_Z_R,`AO12HS_B_R_Z_F);
      (A -=> Z) = (`AO12HS_A_F_Z_R,`AO12HS_A_R_Z_F);

   endspecify
`endif


endmodule // AO12HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:55 and Version :1.1 //
 
//  START 
// CELL AO12NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO12NHS_H_F_Z_F 0.1
`define AO12NHS_H_R_Z_R 0.1
`define AO12NHS_G_F_Z_F 0.1
`define AO12NHS_G_R_Z_R 0.1
`define AO12NHS_F_F_Z_F 0.1
`define AO12NHS_F_R_Z_R 0.1
`define AO12NHS_E_F_Z_F 0.1
`define AO12NHS_E_R_Z_R 0.1
`define AO12NHS_D_F_Z_F 0.1
`define AO12NHS_D_R_Z_R 0.1
`define AO12NHS_C_F_Z_F 0.1
`define AO12NHS_C_R_Z_R 0.1
`define AO12NHS_B_F_Z_F 0.1
`define AO12NHS_B_R_Z_R 0.1
`define AO12NHS_A_F_Z_F 0.1
`define AO12NHS_A_R_Z_R 0.1

module AO12NHS (Z, A, B, C, D, E, F, G, H);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;
   input G;
   input H;


   or  u0 (OrAB_, A, B);
   or  u1 (OrCD_, C, D);
   or  u2 (OrEF_, E, F);
   or  u3 (OrGH_, G, H);
   and  u4 (Z, OrAB_, OrCD_, OrEF_, OrGH_);


`ifdef functional
`else
   specify

      (H +=> Z) = (`AO12NHS_H_R_Z_R,`AO12NHS_H_F_Z_F);
      (G +=> Z) = (`AO12NHS_G_R_Z_R,`AO12NHS_G_F_Z_F);
      (F +=> Z) = (`AO12NHS_F_R_Z_R,`AO12NHS_F_F_Z_F);
      (E +=> Z) = (`AO12NHS_E_R_Z_R,`AO12NHS_E_F_Z_F);
      (D +=> Z) = (`AO12NHS_D_R_Z_R,`AO12NHS_D_F_Z_F);
      (C +=> Z) = (`AO12NHS_C_R_Z_R,`AO12NHS_C_F_Z_F);
      (B +=> Z) = (`AO12NHS_B_R_Z_R,`AO12NHS_B_F_Z_F);
      (A +=> Z) = (`AO12NHS_A_R_Z_R,`AO12NHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO12NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:55 and Version :1.1 //
 
//  START 
// CELL AO12NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO12NHSP_H_F_Z_F 0.1
`define AO12NHSP_H_R_Z_R 0.1
`define AO12NHSP_G_F_Z_F 0.1
`define AO12NHSP_G_R_Z_R 0.1
`define AO12NHSP_F_F_Z_F 0.1
`define AO12NHSP_F_R_Z_R 0.1
`define AO12NHSP_E_F_Z_F 0.1
`define AO12NHSP_E_R_Z_R 0.1
`define AO12NHSP_D_F_Z_F 0.1
`define AO12NHSP_D_R_Z_R 0.1
`define AO12NHSP_C_F_Z_F 0.1
`define AO12NHSP_C_R_Z_R 0.1
`define AO12NHSP_B_F_Z_F 0.1
`define AO12NHSP_B_R_Z_R 0.1
`define AO12NHSP_A_F_Z_F 0.1
`define AO12NHSP_A_R_Z_R 0.1

module AO12NHSP (Z, A, B, C, D, E, F, G, H);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;
   input G;
   input H;


   or  u0 (OrAB_, A, B);
   or  u1 (OrCD_, C, D);
   or  u2 (OrEF_, E, F);
   or  u3 (OrGH_, G, H);
   and  u4 (Z, OrAB_, OrCD_, OrEF_, OrGH_);


`ifdef functional
`else
   specify

      (H +=> Z) = (`AO12NHSP_H_R_Z_R,`AO12NHSP_H_F_Z_F);
      (G +=> Z) = (`AO12NHSP_G_R_Z_R,`AO12NHSP_G_F_Z_F);
      (F +=> Z) = (`AO12NHSP_F_R_Z_R,`AO12NHSP_F_F_Z_F);
      (E +=> Z) = (`AO12NHSP_E_R_Z_R,`AO12NHSP_E_F_Z_F);
      (D +=> Z) = (`AO12NHSP_D_R_Z_R,`AO12NHSP_D_F_Z_F);
      (C +=> Z) = (`AO12NHSP_C_R_Z_R,`AO12NHSP_C_F_Z_F);
      (B +=> Z) = (`AO12NHSP_B_R_Z_R,`AO12NHSP_B_F_Z_F);
      (A +=> Z) = (`AO12NHSP_A_R_Z_R,`AO12NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO12NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:03:55 and Version :1.1 //
 
//  START 
// CELL AO13HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO13HSX05_E_F_Z_R 0.1
`define AO13HSX05_E_R_Z_F 0.1
`define AO13HSX05_D_F_Z_R 0.1
`define AO13HSX05_D_R_Z_F 0.1
`define AO13HSX05_C_F_Z_R 0.1
`define AO13HSX05_C_R_Z_F 0.1
`define AO13HSX05_B_F_Z_R 0.1
`define AO13HSX05_B_R_Z_F 0.1
`define AO13HSX05_A_F_Z_R 0.1
`define AO13HSX05_A_R_Z_F 0.1

module AO13HSX05 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   nand  u0 (Z, OrCDE_, OrABE_);
   or  u1 (OrABE_, A, B, E);
   or  u2 (OrCDE_, C, D, E);


`ifdef functional
`else
   specify

      (E -=> Z) = (`AO13HSX05_E_F_Z_R,`AO13HSX05_E_R_Z_F);
      (D -=> Z) = (`AO13HSX05_D_F_Z_R,`AO13HSX05_D_R_Z_F);
      (C -=> Z) = (`AO13HSX05_C_F_Z_R,`AO13HSX05_C_R_Z_F);
      (B -=> Z) = (`AO13HSX05_B_F_Z_R,`AO13HSX05_B_R_Z_F);
      (A -=> Z) = (`AO13HSX05_A_F_Z_R,`AO13HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // AO13HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:04:13 and Version :1.1 //
 
//  START 
// CELL AO13HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO13HS_E_F_Z_R 0.1
`define AO13HS_E_R_Z_F 0.1
`define AO13HS_D_F_Z_R 0.1
`define AO13HS_D_R_Z_F 0.1
`define AO13HS_C_F_Z_R 0.1
`define AO13HS_C_R_Z_F 0.1
`define AO13HS_B_F_Z_R 0.1
`define AO13HS_B_R_Z_F 0.1
`define AO13HS_A_F_Z_R 0.1
`define AO13HS_A_R_Z_F 0.1

module AO13HS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   nand  u0 (Z, OrCDE_, OrABE_);
   or  u1 (OrABE_, A, B, E);
   or  u2 (OrCDE_, C, D, E);


`ifdef functional
`else
   specify

      (E -=> Z) = (`AO13HS_E_F_Z_R,`AO13HS_E_R_Z_F);
      (D -=> Z) = (`AO13HS_D_F_Z_R,`AO13HS_D_R_Z_F);
      (C -=> Z) = (`AO13HS_C_F_Z_R,`AO13HS_C_R_Z_F);
      (B -=> Z) = (`AO13HS_B_F_Z_R,`AO13HS_B_R_Z_F);
      (A -=> Z) = (`AO13HS_A_F_Z_R,`AO13HS_A_R_Z_F);

   endspecify
`endif


endmodule // AO13HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:04:13 and Version :1.1 //
 
//  START 
// CELL AO13NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO13NHS_E_F_Z_F 0.1
`define AO13NHS_E_R_Z_R 0.1
`define AO13NHS_D_F_Z_F 0.1
`define AO13NHS_D_R_Z_R 0.1
`define AO13NHS_C_F_Z_F 0.1
`define AO13NHS_C_R_Z_R 0.1
`define AO13NHS_B_F_Z_F 0.1
`define AO13NHS_B_R_Z_R 0.1
`define AO13NHS_A_F_Z_F 0.1
`define AO13NHS_A_R_Z_R 0.1

module AO13NHS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   or  u0 (OrCDE_, C, D, E);
   or  u1 (OrABE_, A, B, E);
   and  u2 (Z, OrCDE_, OrABE_);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO13NHS_E_R_Z_R,`AO13NHS_E_F_Z_F);
      (D +=> Z) = (`AO13NHS_D_R_Z_R,`AO13NHS_D_F_Z_F);
      (C +=> Z) = (`AO13NHS_C_R_Z_R,`AO13NHS_C_F_Z_F);
      (B +=> Z) = (`AO13NHS_B_R_Z_R,`AO13NHS_B_F_Z_F);
      (A +=> Z) = (`AO13NHS_A_R_Z_R,`AO13NHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO13NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:04:13 and Version :1.1 //
 
//  START 
// CELL AO13NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO13NHSP_E_F_Z_F 0.1
`define AO13NHSP_E_R_Z_R 0.1
`define AO13NHSP_D_F_Z_F 0.1
`define AO13NHSP_D_R_Z_R 0.1
`define AO13NHSP_C_F_Z_F 0.1
`define AO13NHSP_C_R_Z_R 0.1
`define AO13NHSP_B_F_Z_F 0.1
`define AO13NHSP_B_R_Z_R 0.1
`define AO13NHSP_A_F_Z_F 0.1
`define AO13NHSP_A_R_Z_R 0.1

module AO13NHSP (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   or  u0 (OrCDE_, C, D, E);
   or  u1 (OrABE_, A, B, E);
   and  u2 (Z, OrCDE_, OrABE_);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO13NHSP_E_R_Z_R,`AO13NHSP_E_F_Z_F);
      (D +=> Z) = (`AO13NHSP_D_R_Z_R,`AO13NHSP_D_F_Z_F);
      (C +=> Z) = (`AO13NHSP_C_R_Z_R,`AO13NHSP_C_F_Z_F);
      (B +=> Z) = (`AO13NHSP_B_R_Z_R,`AO13NHSP_B_F_Z_F);
      (A +=> Z) = (`AO13NHSP_A_R_Z_R,`AO13NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO13NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:04:13 and Version :1.1 //
 
//  START 
// CELL AO14HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO14HS_F_F_Z_R 0.1
`define AO14HS_F_R_Z_F 0.1
`define AO14HS_E_F_Z_R 0.1
`define AO14HS_E_R_Z_F 0.1
`define AO14HS_D_F_Z_R 0.1
`define AO14HS_D_R_Z_F 0.1
`define AO14HS_C_F_Z_R 0.1
`define AO14HS_C_R_Z_F 0.1
`define AO14HS_B_F_Z_R 0.1
`define AO14HS_B_R_Z_F 0.1
`define AO14HS_A_F_Z_R 0.1
`define AO14HS_A_R_Z_F 0.1

module AO14HS (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   and  u0 (AndABC_, A, B, C);
   and  u1 (AndDEF_, D, E, F);
   nor  u2 (Z, AndABC_, AndDEF_);


`ifdef functional
`else
   specify

      (F -=> Z) = (`AO14HS_F_F_Z_R,`AO14HS_F_R_Z_F);
      (E -=> Z) = (`AO14HS_E_F_Z_R,`AO14HS_E_R_Z_F);
      (D -=> Z) = (`AO14HS_D_F_Z_R,`AO14HS_D_R_Z_F);
      (C -=> Z) = (`AO14HS_C_F_Z_R,`AO14HS_C_R_Z_F);
      (B -=> Z) = (`AO14HS_B_F_Z_R,`AO14HS_B_R_Z_F);
      (A -=> Z) = (`AO14HS_A_F_Z_R,`AO14HS_A_R_Z_F);

   endspecify
`endif


endmodule // AO14HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:04:26 and Version :1.1 //
 
//  START 
// CELL AO14HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO14HSP_F_F_Z_R 0.1
`define AO14HSP_F_R_Z_F 0.1
`define AO14HSP_E_F_Z_R 0.1
`define AO14HSP_E_R_Z_F 0.1
`define AO14HSP_D_F_Z_R 0.1
`define AO14HSP_D_R_Z_F 0.1
`define AO14HSP_C_F_Z_R 0.1
`define AO14HSP_C_R_Z_F 0.1
`define AO14HSP_B_F_Z_R 0.1
`define AO14HSP_B_R_Z_F 0.1
`define AO14HSP_A_F_Z_R 0.1
`define AO14HSP_A_R_Z_F 0.1

module AO14HSP (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   and  u0 (AndABC_, A, B, C);
   and  u1 (AndDEF_, D, E, F);
   nor  u2 (Z, AndABC_, AndDEF_);


`ifdef functional
`else
   specify

      (F -=> Z) = (`AO14HSP_F_F_Z_R,`AO14HSP_F_R_Z_F);
      (E -=> Z) = (`AO14HSP_E_F_Z_R,`AO14HSP_E_R_Z_F);
      (D -=> Z) = (`AO14HSP_D_F_Z_R,`AO14HSP_D_R_Z_F);
      (C -=> Z) = (`AO14HSP_C_F_Z_R,`AO14HSP_C_R_Z_F);
      (B -=> Z) = (`AO14HSP_B_F_Z_R,`AO14HSP_B_R_Z_F);
      (A -=> Z) = (`AO14HSP_A_F_Z_R,`AO14HSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO14HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:04:26 and Version :1.1 //
 
//  START 
// CELL AO14HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO14HSX4_F_F_Z_R 0.1
`define AO14HSX4_F_R_Z_F 0.1
`define AO14HSX4_E_F_Z_R 0.1
`define AO14HSX4_E_R_Z_F 0.1
`define AO14HSX4_D_F_Z_R 0.1
`define AO14HSX4_D_R_Z_F 0.1
`define AO14HSX4_C_F_Z_R 0.1
`define AO14HSX4_C_R_Z_F 0.1
`define AO14HSX4_B_F_Z_R 0.1
`define AO14HSX4_B_R_Z_F 0.1
`define AO14HSX4_A_F_Z_R 0.1
`define AO14HSX4_A_R_Z_F 0.1

module AO14HSX4 (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   and  u0 (AndABC_, A, B, C);
   and  u1 (AndDEF_, D, E, F);
   nor  u2 (Z, AndABC_, AndDEF_);


`ifdef functional
`else
   specify

      (F -=> Z) = (`AO14HSX4_F_F_Z_R,`AO14HSX4_F_R_Z_F);
      (E -=> Z) = (`AO14HSX4_E_F_Z_R,`AO14HSX4_E_R_Z_F);
      (D -=> Z) = (`AO14HSX4_D_F_Z_R,`AO14HSX4_D_R_Z_F);
      (C -=> Z) = (`AO14HSX4_C_F_Z_R,`AO14HSX4_C_R_Z_F);
      (B -=> Z) = (`AO14HSX4_B_F_Z_R,`AO14HSX4_B_R_Z_F);
      (A -=> Z) = (`AO14HSX4_A_F_Z_R,`AO14HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO14HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:04:26 and Version :1.1 //
 
//  START 
// CELL AO14HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO14HSX8_F_F_Z_R 0.1
`define AO14HSX8_F_R_Z_F 0.1
`define AO14HSX8_E_F_Z_R 0.1
`define AO14HSX8_E_R_Z_F 0.1
`define AO14HSX8_D_F_Z_R 0.1
`define AO14HSX8_D_R_Z_F 0.1
`define AO14HSX8_C_F_Z_R 0.1
`define AO14HSX8_C_R_Z_F 0.1
`define AO14HSX8_B_F_Z_R 0.1
`define AO14HSX8_B_R_Z_F 0.1
`define AO14HSX8_A_F_Z_R 0.1
`define AO14HSX8_A_R_Z_F 0.1

module AO14HSX8 (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   and  u0 (AndABC_, A, B, C);
   and  u1 (AndDEF_, D, E, F);
   nor  u2 (Z, AndABC_, AndDEF_);


`ifdef functional
`else
   specify

      (F -=> Z) = (`AO14HSX8_F_F_Z_R,`AO14HSX8_F_R_Z_F);
      (E -=> Z) = (`AO14HSX8_E_F_Z_R,`AO14HSX8_E_R_Z_F);
      (D -=> Z) = (`AO14HSX8_D_F_Z_R,`AO14HSX8_D_R_Z_F);
      (C -=> Z) = (`AO14HSX8_C_F_Z_R,`AO14HSX8_C_R_Z_F);
      (B -=> Z) = (`AO14HSX8_B_F_Z_R,`AO14HSX8_B_R_Z_F);
      (A -=> Z) = (`AO14HSX8_A_F_Z_R,`AO14HSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AO14HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:04:26 and Version :1.1 //
 
//  START 
// CELL AO14NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO14NHS_F_F_Z_F 0.1
`define AO14NHS_F_R_Z_R 0.1
`define AO14NHS_E_F_Z_F 0.1
`define AO14NHS_E_R_Z_R 0.1
`define AO14NHS_D_F_Z_F 0.1
`define AO14NHS_D_R_Z_R 0.1
`define AO14NHS_C_F_Z_F 0.1
`define AO14NHS_C_R_Z_R 0.1
`define AO14NHS_B_F_Z_F 0.1
`define AO14NHS_B_R_Z_R 0.1
`define AO14NHS_A_F_Z_F 0.1
`define AO14NHS_A_R_Z_R 0.1

module AO14NHS (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   and  u0 (AndABC_, A, B, C);
   and  u1 (AndDEF_, D, E, F);
   or  u2 (Z, AndABC_, AndDEF_);


`ifdef functional
`else
   specify

      (F +=> Z) = (`AO14NHS_F_R_Z_R,`AO14NHS_F_F_Z_F);
      (E +=> Z) = (`AO14NHS_E_R_Z_R,`AO14NHS_E_F_Z_F);
      (D +=> Z) = (`AO14NHS_D_R_Z_R,`AO14NHS_D_F_Z_F);
      (C +=> Z) = (`AO14NHS_C_R_Z_R,`AO14NHS_C_F_Z_F);
      (B +=> Z) = (`AO14NHS_B_R_Z_R,`AO14NHS_B_F_Z_F);
      (A +=> Z) = (`AO14NHS_A_R_Z_R,`AO14NHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO14NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:04:26 and Version :1.1 //
 
//  START 
// CELL AO14NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO14NHSP_F_F_Z_F 0.1
`define AO14NHSP_F_R_Z_R 0.1
`define AO14NHSP_E_F_Z_F 0.1
`define AO14NHSP_E_R_Z_R 0.1
`define AO14NHSP_D_F_Z_F 0.1
`define AO14NHSP_D_R_Z_R 0.1
`define AO14NHSP_C_F_Z_F 0.1
`define AO14NHSP_C_R_Z_R 0.1
`define AO14NHSP_B_F_Z_F 0.1
`define AO14NHSP_B_R_Z_R 0.1
`define AO14NHSP_A_F_Z_F 0.1
`define AO14NHSP_A_R_Z_R 0.1

module AO14NHSP (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   and  u0 (AndABC_, A, B, C);
   and  u1 (AndDEF_, D, E, F);
   or  u2 (Z, AndABC_, AndDEF_);


`ifdef functional
`else
   specify

      (F +=> Z) = (`AO14NHSP_F_R_Z_R,`AO14NHSP_F_F_Z_F);
      (E +=> Z) = (`AO14NHSP_E_R_Z_R,`AO14NHSP_E_F_Z_F);
      (D +=> Z) = (`AO14NHSP_D_R_Z_R,`AO14NHSP_D_F_Z_F);
      (C +=> Z) = (`AO14NHSP_C_R_Z_R,`AO14NHSP_C_F_Z_F);
      (B +=> Z) = (`AO14NHSP_B_R_Z_R,`AO14NHSP_B_F_Z_F);
      (A +=> Z) = (`AO14NHSP_A_R_Z_R,`AO14NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO14NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:04:26 and Version :1.1 //
 
//  START 
// CELL AO14NHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO14NHSX4_F_F_Z_F 0.1
`define AO14NHSX4_F_R_Z_R 0.1
`define AO14NHSX4_E_F_Z_F 0.1
`define AO14NHSX4_E_R_Z_R 0.1
`define AO14NHSX4_D_F_Z_F 0.1
`define AO14NHSX4_D_R_Z_R 0.1
`define AO14NHSX4_C_F_Z_F 0.1
`define AO14NHSX4_C_R_Z_R 0.1
`define AO14NHSX4_B_F_Z_F 0.1
`define AO14NHSX4_B_R_Z_R 0.1
`define AO14NHSX4_A_F_Z_F 0.1
`define AO14NHSX4_A_R_Z_R 0.1

module AO14NHSX4 (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   and  u0 (AndABC_, A, B, C);
   and  u1 (AndDEF_, D, E, F);
   or  u2 (Z, AndABC_, AndDEF_);


`ifdef functional
`else
   specify

      (F +=> Z) = (`AO14NHSX4_F_R_Z_R,`AO14NHSX4_F_F_Z_F);
      (E +=> Z) = (`AO14NHSX4_E_R_Z_R,`AO14NHSX4_E_F_Z_F);
      (D +=> Z) = (`AO14NHSX4_D_R_Z_R,`AO14NHSX4_D_F_Z_F);
      (C +=> Z) = (`AO14NHSX4_C_R_Z_R,`AO14NHSX4_C_F_Z_F);
      (B +=> Z) = (`AO14NHSX4_B_R_Z_R,`AO14NHSX4_B_F_Z_F);
      (A +=> Z) = (`AO14NHSX4_A_R_Z_R,`AO14NHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO14NHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:04:26 and Version :1.1 //
 
//  START 
// CELL AO14NHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO14NHSX8_F_F_Z_F 0.1
`define AO14NHSX8_F_R_Z_R 0.1
`define AO14NHSX8_E_F_Z_F 0.1
`define AO14NHSX8_E_R_Z_R 0.1
`define AO14NHSX8_D_F_Z_F 0.1
`define AO14NHSX8_D_R_Z_R 0.1
`define AO14NHSX8_C_F_Z_F 0.1
`define AO14NHSX8_C_R_Z_R 0.1
`define AO14NHSX8_B_F_Z_F 0.1
`define AO14NHSX8_B_R_Z_R 0.1
`define AO14NHSX8_A_F_Z_F 0.1
`define AO14NHSX8_A_R_Z_R 0.1

module AO14NHSX8 (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   and  u0 (AndABC_, A, B, C);
   and  u1 (AndDEF_, D, E, F);
   or  u2 (Z, AndABC_, AndDEF_);


`ifdef functional
`else
   specify

      (F +=> Z) = (`AO14NHSX8_F_R_Z_R,`AO14NHSX8_F_F_Z_F);
      (E +=> Z) = (`AO14NHSX8_E_R_Z_R,`AO14NHSX8_E_F_Z_F);
      (D +=> Z) = (`AO14NHSX8_D_R_Z_R,`AO14NHSX8_D_F_Z_F);
      (C +=> Z) = (`AO14NHSX8_C_R_Z_R,`AO14NHSX8_C_F_Z_F);
      (B +=> Z) = (`AO14NHSX8_B_R_Z_R,`AO14NHSX8_B_F_Z_F);
      (A +=> Z) = (`AO14NHSX8_A_R_Z_R,`AO14NHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO14NHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:04:26 and Version :1.1 //
 
//  START 
// CELL AO15HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO15HSX05_F_F_Z_R 0.1
`define AO15HSX05_F_R_Z_F 0.1
`define AO15HSX05_E_F_Z_R 0.1
`define AO15HSX05_E_R_Z_F 0.1
`define AO15HSX05_D_F_Z_R 0.1
`define AO15HSX05_D_R_Z_F 0.1
`define AO15HSX05_C_F_Z_R 0.1
`define AO15HSX05_C_R_Z_F 0.1
`define AO15HSX05_B_F_Z_R 0.1
`define AO15HSX05_B_R_Z_F 0.1
`define AO15HSX05_A_F_Z_R 0.1
`define AO15HSX05_A_R_Z_F 0.1

module AO15HSX05 (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   nand  u0 (Z, OrABC_, OrDEF_);
   or  u1 (OrDEF_, D, E, F);
   or  u2 (OrABC_, A, B, C);


`ifdef functional
`else
   specify

      (F -=> Z) = (`AO15HSX05_F_F_Z_R,`AO15HSX05_F_R_Z_F);
      (E -=> Z) = (`AO15HSX05_E_F_Z_R,`AO15HSX05_E_R_Z_F);
      (D -=> Z) = (`AO15HSX05_D_F_Z_R,`AO15HSX05_D_R_Z_F);
      (C -=> Z) = (`AO15HSX05_C_F_Z_R,`AO15HSX05_C_R_Z_F);
      (B -=> Z) = (`AO15HSX05_B_F_Z_R,`AO15HSX05_B_R_Z_F);
      (A -=> Z) = (`AO15HSX05_A_F_Z_R,`AO15HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // AO15HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:04:38 and Version :1.1 //
 
//  START 
// CELL AO15HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO15HS_F_F_Z_R 0.1
`define AO15HS_F_R_Z_F 0.1
`define AO15HS_E_F_Z_R 0.1
`define AO15HS_E_R_Z_F 0.1
`define AO15HS_D_F_Z_R 0.1
`define AO15HS_D_R_Z_F 0.1
`define AO15HS_C_F_Z_R 0.1
`define AO15HS_C_R_Z_F 0.1
`define AO15HS_B_F_Z_R 0.1
`define AO15HS_B_R_Z_F 0.1
`define AO15HS_A_F_Z_R 0.1
`define AO15HS_A_R_Z_F 0.1

module AO15HS (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   nand  u0 (Z, OrABC_, OrDEF_);
   or  u1 (OrDEF_, D, E, F);
   or  u2 (OrABC_, A, B, C);


`ifdef functional
`else
   specify

      (F -=> Z) = (`AO15HS_F_F_Z_R,`AO15HS_F_R_Z_F);
      (E -=> Z) = (`AO15HS_E_F_Z_R,`AO15HS_E_R_Z_F);
      (D -=> Z) = (`AO15HS_D_F_Z_R,`AO15HS_D_R_Z_F);
      (C -=> Z) = (`AO15HS_C_F_Z_R,`AO15HS_C_R_Z_F);
      (B -=> Z) = (`AO15HS_B_F_Z_R,`AO15HS_B_R_Z_F);
      (A -=> Z) = (`AO15HS_A_F_Z_R,`AO15HS_A_R_Z_F);

   endspecify
`endif


endmodule // AO15HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:04:38 and Version :1.1 //
 
//  START 
// CELL AO15NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO15NHS_F_F_Z_F 0.1
`define AO15NHS_F_R_Z_R 0.1
`define AO15NHS_E_F_Z_F 0.1
`define AO15NHS_E_R_Z_R 0.1
`define AO15NHS_D_F_Z_F 0.1
`define AO15NHS_D_R_Z_R 0.1
`define AO15NHS_C_F_Z_F 0.1
`define AO15NHS_C_R_Z_R 0.1
`define AO15NHS_B_F_Z_F 0.1
`define AO15NHS_B_R_Z_R 0.1
`define AO15NHS_A_F_Z_F 0.1
`define AO15NHS_A_R_Z_R 0.1

module AO15NHS (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   or  u0 (OrABC_, A, B, C);
   or  u1 (OrDEF_, D, E, F);
   and  u2 (Z, OrABC_, OrDEF_);


`ifdef functional
`else
   specify

      (F +=> Z) = (`AO15NHS_F_R_Z_R,`AO15NHS_F_F_Z_F);
      (E +=> Z) = (`AO15NHS_E_R_Z_R,`AO15NHS_E_F_Z_F);
      (D +=> Z) = (`AO15NHS_D_R_Z_R,`AO15NHS_D_F_Z_F);
      (C +=> Z) = (`AO15NHS_C_R_Z_R,`AO15NHS_C_F_Z_F);
      (B +=> Z) = (`AO15NHS_B_R_Z_R,`AO15NHS_B_F_Z_F);
      (A +=> Z) = (`AO15NHS_A_R_Z_R,`AO15NHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO15NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:04:38 and Version :1.1 //
 
//  START 
// CELL AO15NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO15NHSP_F_F_Z_F 0.1
`define AO15NHSP_F_R_Z_R 0.1
`define AO15NHSP_E_F_Z_F 0.1
`define AO15NHSP_E_R_Z_R 0.1
`define AO15NHSP_D_F_Z_F 0.1
`define AO15NHSP_D_R_Z_R 0.1
`define AO15NHSP_C_F_Z_F 0.1
`define AO15NHSP_C_R_Z_R 0.1
`define AO15NHSP_B_F_Z_F 0.1
`define AO15NHSP_B_R_Z_R 0.1
`define AO15NHSP_A_F_Z_F 0.1
`define AO15NHSP_A_R_Z_R 0.1

module AO15NHSP (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   or  u0 (OrABC_, A, B, C);
   or  u1 (OrDEF_, D, E, F);
   and  u2 (Z, OrABC_, OrDEF_);


`ifdef functional
`else
   specify

      (F +=> Z) = (`AO15NHSP_F_R_Z_R,`AO15NHSP_F_F_Z_F);
      (E +=> Z) = (`AO15NHSP_E_R_Z_R,`AO15NHSP_E_F_Z_F);
      (D +=> Z) = (`AO15NHSP_D_R_Z_R,`AO15NHSP_D_F_Z_F);
      (C +=> Z) = (`AO15NHSP_C_R_Z_R,`AO15NHSP_C_F_Z_F);
      (B +=> Z) = (`AO15NHSP_B_R_Z_R,`AO15NHSP_B_F_Z_F);
      (A +=> Z) = (`AO15NHSP_A_R_Z_R,`AO15NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO15NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:04:38 and Version :1.1 //
 
//  START 
// CELL AO16HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO16HS_H_F_Z_R 0.1
`define AO16HS_H_R_Z_F 0.1
`define AO16HS_G_F_Z_R 0.1
`define AO16HS_G_R_Z_F 0.1
`define AO16HS_F_F_Z_R 0.1
`define AO16HS_F_R_Z_F 0.1
`define AO16HS_E_F_Z_R 0.1
`define AO16HS_E_R_Z_F 0.1
`define AO16HS_D_F_Z_R 0.1
`define AO16HS_D_R_Z_F 0.1
`define AO16HS_C_F_Z_R 0.1
`define AO16HS_C_R_Z_F 0.1
`define AO16HS_B_F_Z_R 0.1
`define AO16HS_B_R_Z_F 0.1
`define AO16HS_A_F_Z_R 0.1
`define AO16HS_A_R_Z_F 0.1

module AO16HS (Z, A, B, C, D, E, F, G, H);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;
   input G;
   input H;


   and  u0 (AndABCD_, A, B, C, D);
   and  u1 (AndEFGH_, E, F, G, H);
   nor  u2 (Z, AndABCD_, AndEFGH_);


`ifdef functional
`else
   specify

      (H -=> Z) = (`AO16HS_H_F_Z_R,`AO16HS_H_R_Z_F);
      (G -=> Z) = (`AO16HS_G_F_Z_R,`AO16HS_G_R_Z_F);
      (F -=> Z) = (`AO16HS_F_F_Z_R,`AO16HS_F_R_Z_F);
      (E -=> Z) = (`AO16HS_E_F_Z_R,`AO16HS_E_R_Z_F);
      (D -=> Z) = (`AO16HS_D_F_Z_R,`AO16HS_D_R_Z_F);
      (C -=> Z) = (`AO16HS_C_F_Z_R,`AO16HS_C_R_Z_F);
      (B -=> Z) = (`AO16HS_B_F_Z_R,`AO16HS_B_R_Z_F);
      (A -=> Z) = (`AO16HS_A_F_Z_R,`AO16HS_A_R_Z_F);

   endspecify
`endif


endmodule // AO16HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:04:50 and Version :1.1 //
 
//  START 
// CELL AO16NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO16NHS_H_F_Z_F 0.1
`define AO16NHS_H_R_Z_R 0.1
`define AO16NHS_G_F_Z_F 0.1
`define AO16NHS_G_R_Z_R 0.1
`define AO16NHS_F_F_Z_F 0.1
`define AO16NHS_F_R_Z_R 0.1
`define AO16NHS_E_F_Z_F 0.1
`define AO16NHS_E_R_Z_R 0.1
`define AO16NHS_D_F_Z_F 0.1
`define AO16NHS_D_R_Z_R 0.1
`define AO16NHS_C_F_Z_F 0.1
`define AO16NHS_C_R_Z_R 0.1
`define AO16NHS_B_F_Z_F 0.1
`define AO16NHS_B_R_Z_R 0.1
`define AO16NHS_A_F_Z_F 0.1
`define AO16NHS_A_R_Z_R 0.1

module AO16NHS (Z, A, B, C, D, E, F, G, H);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;
   input G;
   input H;


   and  u0 (AndABCD_, A, B, C, D);
   and  u1 (AndEFGH_, E, F, G, H);
   or  u2 (Z, AndABCD_, AndEFGH_);


`ifdef functional
`else
   specify

      (H +=> Z) = (`AO16NHS_H_R_Z_R,`AO16NHS_H_F_Z_F);
      (G +=> Z) = (`AO16NHS_G_R_Z_R,`AO16NHS_G_F_Z_F);
      (F +=> Z) = (`AO16NHS_F_R_Z_R,`AO16NHS_F_F_Z_F);
      (E +=> Z) = (`AO16NHS_E_R_Z_R,`AO16NHS_E_F_Z_F);
      (D +=> Z) = (`AO16NHS_D_R_Z_R,`AO16NHS_D_F_Z_F);
      (C +=> Z) = (`AO16NHS_C_R_Z_R,`AO16NHS_C_F_Z_F);
      (B +=> Z) = (`AO16NHS_B_R_Z_R,`AO16NHS_B_F_Z_F);
      (A +=> Z) = (`AO16NHS_A_R_Z_R,`AO16NHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO16NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:04:50 and Version :1.1 //
 
//  START 
// CELL AO16NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO16NHSP_H_F_Z_F 0.1
`define AO16NHSP_H_R_Z_R 0.1
`define AO16NHSP_G_F_Z_F 0.1
`define AO16NHSP_G_R_Z_R 0.1
`define AO16NHSP_F_F_Z_F 0.1
`define AO16NHSP_F_R_Z_R 0.1
`define AO16NHSP_E_F_Z_F 0.1
`define AO16NHSP_E_R_Z_R 0.1
`define AO16NHSP_D_F_Z_F 0.1
`define AO16NHSP_D_R_Z_R 0.1
`define AO16NHSP_C_F_Z_F 0.1
`define AO16NHSP_C_R_Z_R 0.1
`define AO16NHSP_B_F_Z_F 0.1
`define AO16NHSP_B_R_Z_R 0.1
`define AO16NHSP_A_F_Z_F 0.1
`define AO16NHSP_A_R_Z_R 0.1

module AO16NHSP (Z, A, B, C, D, E, F, G, H);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;
   input G;
   input H;


   and  u0 (AndABCD_, A, B, C, D);
   and  u1 (AndEFGH_, E, F, G, H);
   or  u2 (Z, AndABCD_, AndEFGH_);


`ifdef functional
`else
   specify

      (H +=> Z) = (`AO16NHSP_H_R_Z_R,`AO16NHSP_H_F_Z_F);
      (G +=> Z) = (`AO16NHSP_G_R_Z_R,`AO16NHSP_G_F_Z_F);
      (F +=> Z) = (`AO16NHSP_F_R_Z_R,`AO16NHSP_F_F_Z_F);
      (E +=> Z) = (`AO16NHSP_E_R_Z_R,`AO16NHSP_E_F_Z_F);
      (D +=> Z) = (`AO16NHSP_D_R_Z_R,`AO16NHSP_D_F_Z_F);
      (C +=> Z) = (`AO16NHSP_C_R_Z_R,`AO16NHSP_C_F_Z_F);
      (B +=> Z) = (`AO16NHSP_B_R_Z_R,`AO16NHSP_B_F_Z_F);
      (A +=> Z) = (`AO16NHSP_A_R_Z_R,`AO16NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO16NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:04:50 and Version :1.1 //
 
//  START 
// CELL AO17HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO17HSX05_D_F_Z_R 0.1
`define AO17HSX05_D_R_Z_F 0.1
`define AO17HSX05_C_F_Z_R 0.1
`define AO17HSX05_C_R_Z_F 0.1
`define AO17HSX05_B_F_Z_R 0.1
`define AO17HSX05_B_R_Z_F 0.1
`define AO17HSX05_A_F_Z_R 0.1
`define AO17HSX05_A_R_Z_F 0.1

module AO17HSX05 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (AndAB_, A, B);
   or  u1 (OrAndAB_C_, AndAB_, C);
   nand  u2 (Z, OrAndAB_C_, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO17HSX05_D_F_Z_R,`AO17HSX05_D_R_Z_F);
      (C -=> Z) = (`AO17HSX05_C_F_Z_R,`AO17HSX05_C_R_Z_F);
      (B -=> Z) = (`AO17HSX05_B_F_Z_R,`AO17HSX05_B_R_Z_F);
      (A -=> Z) = (`AO17HSX05_A_F_Z_R,`AO17HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // AO17HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:13 and Version :1.1 //
 
//  START 
// CELL AO17HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO17HS_D_F_Z_R 0.1
`define AO17HS_D_R_Z_F 0.1
`define AO17HS_C_F_Z_R 0.1
`define AO17HS_C_R_Z_F 0.1
`define AO17HS_B_F_Z_R 0.1
`define AO17HS_B_R_Z_F 0.1
`define AO17HS_A_F_Z_R 0.1
`define AO17HS_A_R_Z_F 0.1

module AO17HS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (AndAB_, A, B);
   or  u1 (OrAndAB_C_, AndAB_, C);
   nand  u2 (Z, OrAndAB_C_, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO17HS_D_F_Z_R,`AO17HS_D_R_Z_F);
      (C -=> Z) = (`AO17HS_C_F_Z_R,`AO17HS_C_R_Z_F);
      (B -=> Z) = (`AO17HS_B_F_Z_R,`AO17HS_B_R_Z_F);
      (A -=> Z) = (`AO17HS_A_F_Z_R,`AO17HS_A_R_Z_F);

   endspecify
`endif


endmodule // AO17HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:13 and Version :1.1 //
 
//  START 
// CELL AO17HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO17HSP_D_F_Z_R 0.1
`define AO17HSP_D_R_Z_F 0.1
`define AO17HSP_C_F_Z_R 0.1
`define AO17HSP_C_R_Z_F 0.1
`define AO17HSP_B_F_Z_R 0.1
`define AO17HSP_B_R_Z_F 0.1
`define AO17HSP_A_F_Z_R 0.1
`define AO17HSP_A_R_Z_F 0.1

module AO17HSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (AndAB_, A, B);
   or  u1 (OrAndAB_C_, AndAB_, C);
   nand  u2 (Z, OrAndAB_C_, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO17HSP_D_F_Z_R,`AO17HSP_D_R_Z_F);
      (C -=> Z) = (`AO17HSP_C_F_Z_R,`AO17HSP_C_R_Z_F);
      (B -=> Z) = (`AO17HSP_B_F_Z_R,`AO17HSP_B_R_Z_F);
      (A -=> Z) = (`AO17HSP_A_F_Z_R,`AO17HSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO17HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:13 and Version :1.1 //
 
//  START 
// CELL AO17HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO17HSX4_D_F_Z_R 0.1
`define AO17HSX4_D_R_Z_F 0.1
`define AO17HSX4_C_F_Z_R 0.1
`define AO17HSX4_C_R_Z_F 0.1
`define AO17HSX4_B_F_Z_R 0.1
`define AO17HSX4_B_R_Z_F 0.1
`define AO17HSX4_A_F_Z_R 0.1
`define AO17HSX4_A_R_Z_F 0.1

module AO17HSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (AndAB_, A, B);
   or  u1 (OrAndAB_C_, AndAB_, C);
   nand  u2 (Z, OrAndAB_C_, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO17HSX4_D_F_Z_R,`AO17HSX4_D_R_Z_F);
      (C -=> Z) = (`AO17HSX4_C_F_Z_R,`AO17HSX4_C_R_Z_F);
      (B -=> Z) = (`AO17HSX4_B_F_Z_R,`AO17HSX4_B_R_Z_F);
      (A -=> Z) = (`AO17HSX4_A_F_Z_R,`AO17HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO17HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:13 and Version :1.1 //
 
//  START 
// CELL AO17NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO17NHS_D_F_Z_F 0.1
`define AO17NHS_D_R_Z_R 0.1
`define AO17NHS_C_F_Z_F 0.1
`define AO17NHS_C_R_Z_R 0.1
`define AO17NHS_B_F_Z_F 0.1
`define AO17NHS_B_R_Z_R 0.1
`define AO17NHS_A_F_Z_F 0.1
`define AO17NHS_A_R_Z_R 0.1

module AO17NHS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (AndAB_, A, B);
   or  u1 (OrAndAB_C_, AndAB_, C);
   and  u2 (Z, OrAndAB_C_, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO17NHS_D_R_Z_R,`AO17NHS_D_F_Z_F);
      (C +=> Z) = (`AO17NHS_C_R_Z_R,`AO17NHS_C_F_Z_F);
      (B +=> Z) = (`AO17NHS_B_R_Z_R,`AO17NHS_B_F_Z_F);
      (A +=> Z) = (`AO17NHS_A_R_Z_R,`AO17NHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO17NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:13 and Version :1.1 //
 
//  START 
// CELL AO17NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO17NHSP_D_F_Z_F 0.1
`define AO17NHSP_D_R_Z_R 0.1
`define AO17NHSP_C_F_Z_F 0.1
`define AO17NHSP_C_R_Z_R 0.1
`define AO17NHSP_B_F_Z_F 0.1
`define AO17NHSP_B_R_Z_R 0.1
`define AO17NHSP_A_F_Z_F 0.1
`define AO17NHSP_A_R_Z_R 0.1

module AO17NHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (AndAB_, A, B);
   or  u1 (OrAndAB_C_, AndAB_, C);
   and  u2 (Z, OrAndAB_C_, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO17NHSP_D_R_Z_R,`AO17NHSP_D_F_Z_F);
      (C +=> Z) = (`AO17NHSP_C_R_Z_R,`AO17NHSP_C_F_Z_F);
      (B +=> Z) = (`AO17NHSP_B_R_Z_R,`AO17NHSP_B_F_Z_F);
      (A +=> Z) = (`AO17NHSP_A_R_Z_R,`AO17NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO17NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:13 and Version :1.1 //
 
//  START 
// CELL AO18HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO18HSX05_E_F_Z_R 0.1
`define AO18HSX05_E_R_Z_F 0.1
`define AO18HSX05_D_F_Z_R 0.1
`define AO18HSX05_D_R_Z_F 0.1
`define AO18HSX05_C_F_Z_R 0.1
`define AO18HSX05_C_R_Z_F 0.1
`define AO18HSX05_B_F_Z_R 0.1
`define AO18HSX05_B_R_Z_F 0.1
`define AO18HSX05_A_F_Z_R 0.1
`define AO18HSX05_A_R_Z_F 0.1

module AO18HSX05 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   nor  u0 (Z, AndABE_, AndCDE_);
   and  u1 (AndCDE_, C, D, E);
   and  u2 (AndABE_, A, B, E);


`ifdef functional
`else
   specify

      (E -=> Z) = (`AO18HSX05_E_F_Z_R,`AO18HSX05_E_R_Z_F);
      (D -=> Z) = (`AO18HSX05_D_F_Z_R,`AO18HSX05_D_R_Z_F);
      (C -=> Z) = (`AO18HSX05_C_F_Z_R,`AO18HSX05_C_R_Z_F);
      (B -=> Z) = (`AO18HSX05_B_F_Z_R,`AO18HSX05_B_R_Z_F);
      (A -=> Z) = (`AO18HSX05_A_F_Z_R,`AO18HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // AO18HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:33 and Version :1.1 //
 
//  START 
// CELL AO18HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO18HS_E_F_Z_R 0.1
`define AO18HS_E_R_Z_F 0.1
`define AO18HS_D_F_Z_R 0.1
`define AO18HS_D_R_Z_F 0.1
`define AO18HS_C_F_Z_R 0.1
`define AO18HS_C_R_Z_F 0.1
`define AO18HS_B_F_Z_R 0.1
`define AO18HS_B_R_Z_F 0.1
`define AO18HS_A_F_Z_R 0.1
`define AO18HS_A_R_Z_F 0.1

module AO18HS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   nor  u0 (Z, AndABE_, AndCDE_);
   and  u1 (AndCDE_, C, D, E);
   and  u2 (AndABE_, A, B, E);


`ifdef functional
`else
   specify

      (E -=> Z) = (`AO18HS_E_F_Z_R,`AO18HS_E_R_Z_F);
      (D -=> Z) = (`AO18HS_D_F_Z_R,`AO18HS_D_R_Z_F);
      (C -=> Z) = (`AO18HS_C_F_Z_R,`AO18HS_C_R_Z_F);
      (B -=> Z) = (`AO18HS_B_F_Z_R,`AO18HS_B_R_Z_F);
      (A -=> Z) = (`AO18HS_A_F_Z_R,`AO18HS_A_R_Z_F);

   endspecify
`endif


endmodule // AO18HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:33 and Version :1.1 //
 
//  START 
// CELL AO18NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO18NHS_E_F_Z_F 0.1
`define AO18NHS_E_R_Z_R 0.1
`define AO18NHS_D_F_Z_F 0.1
`define AO18NHS_D_R_Z_R 0.1
`define AO18NHS_C_F_Z_F 0.1
`define AO18NHS_C_R_Z_R 0.1
`define AO18NHS_B_F_Z_F 0.1
`define AO18NHS_B_R_Z_R 0.1
`define AO18NHS_A_F_Z_F 0.1
`define AO18NHS_A_R_Z_R 0.1

module AO18NHS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndABE_, A, B, E);
   and  u1 (AndCDE_, C, D, E);
   or  u2 (Z, AndABE_, AndCDE_);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO18NHS_E_R_Z_R,`AO18NHS_E_F_Z_F);
      (D +=> Z) = (`AO18NHS_D_R_Z_R,`AO18NHS_D_F_Z_F);
      (C +=> Z) = (`AO18NHS_C_R_Z_R,`AO18NHS_C_F_Z_F);
      (B +=> Z) = (`AO18NHS_B_R_Z_R,`AO18NHS_B_F_Z_F);
      (A +=> Z) = (`AO18NHS_A_R_Z_R,`AO18NHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO18NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:33 and Version :1.1 //
 
//  START 
// CELL AO18NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO18NHSP_E_F_Z_F 0.1
`define AO18NHSP_E_R_Z_R 0.1
`define AO18NHSP_D_F_Z_F 0.1
`define AO18NHSP_D_R_Z_R 0.1
`define AO18NHSP_C_F_Z_F 0.1
`define AO18NHSP_C_R_Z_R 0.1
`define AO18NHSP_B_F_Z_F 0.1
`define AO18NHSP_B_R_Z_R 0.1
`define AO18NHSP_A_F_Z_F 0.1
`define AO18NHSP_A_R_Z_R 0.1

module AO18NHSP (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndABE_, A, B, E);
   and  u1 (AndCDE_, C, D, E);
   or  u2 (Z, AndABE_, AndCDE_);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO18NHSP_E_R_Z_R,`AO18NHSP_E_F_Z_F);
      (D +=> Z) = (`AO18NHSP_D_R_Z_R,`AO18NHSP_D_F_Z_F);
      (C +=> Z) = (`AO18NHSP_C_R_Z_R,`AO18NHSP_C_F_Z_F);
      (B +=> Z) = (`AO18NHSP_B_R_Z_R,`AO18NHSP_B_F_Z_F);
      (A +=> Z) = (`AO18NHSP_A_R_Z_R,`AO18NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO18NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:33 and Version :1.1 //
 
//  START 
// CELL AO1AHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1AHS_D_F_Z_R 0.1
`define AO1AHS_D_R_Z_F 0.1
`define AO1AHS_C_F_Z_R 0.1
`define AO1AHS_C_R_Z_F 0.1
`define AO1AHS_B_F_Z_R 0.1
`define AO1AHS_B_R_Z_F 0.1
`define AO1AHS_A_F_Z_F 0.1
`define AO1AHS_A_R_Z_R 0.1

module AO1AHS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAXB_, C, D);
   and  u1 (AndAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO1AHS_D_F_Z_R,`AO1AHS_D_R_Z_F);
      (C -=> Z) = (`AO1AHS_C_F_Z_R,`AO1AHS_C_R_Z_F);
      (B -=> Z) = (`AO1AHS_B_F_Z_R,`AO1AHS_B_R_Z_F);
      (A +=> Z) = (`AO1AHS_A_R_Z_R,`AO1AHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO1AHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:39 and Version :1.1 //
 
//  START 
// CELL AO1AHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1AHSP_D_F_Z_R 0.1
`define AO1AHSP_D_R_Z_F 0.1
`define AO1AHSP_C_F_Z_R 0.1
`define AO1AHSP_C_R_Z_F 0.1
`define AO1AHSP_B_F_Z_R 0.1
`define AO1AHSP_B_R_Z_F 0.1
`define AO1AHSP_A_F_Z_F 0.1
`define AO1AHSP_A_R_Z_R 0.1

module AO1AHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAXB_, C, D);
   and  u1 (AndAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO1AHSP_D_F_Z_R,`AO1AHSP_D_R_Z_F);
      (C -=> Z) = (`AO1AHSP_C_F_Z_R,`AO1AHSP_C_R_Z_F);
      (B -=> Z) = (`AO1AHSP_B_F_Z_R,`AO1AHSP_B_R_Z_F);
      (A +=> Z) = (`AO1AHSP_A_R_Z_R,`AO1AHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO1AHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:39 and Version :1.1 //
 
//  START 
// CELL AO1AHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1AHSX4_D_F_Z_R 0.1
`define AO1AHSX4_D_R_Z_F 0.1
`define AO1AHSX4_C_F_Z_R 0.1
`define AO1AHSX4_C_R_Z_F 0.1
`define AO1AHSX4_B_F_Z_R 0.1
`define AO1AHSX4_B_R_Z_F 0.1
`define AO1AHSX4_A_F_Z_F 0.1
`define AO1AHSX4_A_R_Z_R 0.1

module AO1AHSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAXB_, C, D);
   and  u1 (AndAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO1AHSX4_D_F_Z_R,`AO1AHSX4_D_R_Z_F);
      (C -=> Z) = (`AO1AHSX4_C_F_Z_R,`AO1AHSX4_C_R_Z_F);
      (B -=> Z) = (`AO1AHSX4_B_F_Z_R,`AO1AHSX4_B_R_Z_F);
      (A +=> Z) = (`AO1AHSX4_A_R_Z_R,`AO1AHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO1AHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:39 and Version :1.1 //
 
//  START 
// CELL AO1AHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1AHSX8_D_F_Z_R 0.1
`define AO1AHSX8_D_R_Z_F 0.1
`define AO1AHSX8_C_F_Z_R 0.1
`define AO1AHSX8_C_R_Z_F 0.1
`define AO1AHSX8_B_F_Z_R 0.1
`define AO1AHSX8_B_R_Z_F 0.1
`define AO1AHSX8_A_F_Z_F 0.1
`define AO1AHSX8_A_R_Z_R 0.1

module AO1AHSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAXB_, C, D);
   and  u1 (AndAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO1AHSX8_D_F_Z_R,`AO1AHSX8_D_R_Z_F);
      (C -=> Z) = (`AO1AHSX8_C_F_Z_R,`AO1AHSX8_C_R_Z_F);
      (B -=> Z) = (`AO1AHSX8_B_F_Z_R,`AO1AHSX8_B_R_Z_F);
      (A +=> Z) = (`AO1AHSX8_A_R_Z_R,`AO1AHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO1AHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:39 and Version :1.1 //
 
//  START 
// CELL AO1ANHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1ANHS_D_F_Z_F 0.1
`define AO1ANHS_D_R_Z_R 0.1
`define AO1ANHS_C_F_Z_F 0.1
`define AO1ANHS_C_R_Z_R 0.1
`define AO1ANHS_B_F_Z_F 0.1
`define AO1ANHS_B_R_Z_R 0.1
`define AO1ANHS_A_F_Z_R 0.1
`define AO1ANHS_A_R_Z_F 0.1

module AO1ANHS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, AndAXB_, C, D);
   and  u1 (AndAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO1ANHS_D_R_Z_R,`AO1ANHS_D_F_Z_F);
      (C +=> Z) = (`AO1ANHS_C_R_Z_R,`AO1ANHS_C_F_Z_F);
      (B +=> Z) = (`AO1ANHS_B_R_Z_R,`AO1ANHS_B_F_Z_F);
      (A -=> Z) = (`AO1ANHS_A_F_Z_R,`AO1ANHS_A_R_Z_F);

   endspecify
`endif


endmodule // AO1ANHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:39 and Version :1.1 //
 
//  START 
// CELL AO1ANHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1ANHSP_D_F_Z_F 0.1
`define AO1ANHSP_D_R_Z_R 0.1
`define AO1ANHSP_C_F_Z_F 0.1
`define AO1ANHSP_C_R_Z_R 0.1
`define AO1ANHSP_B_F_Z_F 0.1
`define AO1ANHSP_B_R_Z_R 0.1
`define AO1ANHSP_A_F_Z_R 0.1
`define AO1ANHSP_A_R_Z_F 0.1

module AO1ANHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, AndAXB_, C, D);
   and  u1 (AndAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO1ANHSP_D_R_Z_R,`AO1ANHSP_D_F_Z_F);
      (C +=> Z) = (`AO1ANHSP_C_R_Z_R,`AO1ANHSP_C_F_Z_F);
      (B +=> Z) = (`AO1ANHSP_B_R_Z_R,`AO1ANHSP_B_F_Z_F);
      (A -=> Z) = (`AO1ANHSP_A_F_Z_R,`AO1ANHSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO1ANHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:39 and Version :1.1 //
 
//  START 
// CELL AO1ANHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1ANHSX4_D_F_Z_F 0.1
`define AO1ANHSX4_D_R_Z_R 0.1
`define AO1ANHSX4_C_F_Z_F 0.1
`define AO1ANHSX4_C_R_Z_R 0.1
`define AO1ANHSX4_B_F_Z_F 0.1
`define AO1ANHSX4_B_R_Z_R 0.1
`define AO1ANHSX4_A_F_Z_R 0.1
`define AO1ANHSX4_A_R_Z_F 0.1

module AO1ANHSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, AndAXB_, C, D);
   and  u1 (AndAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO1ANHSX4_D_R_Z_R,`AO1ANHSX4_D_F_Z_F);
      (C +=> Z) = (`AO1ANHSX4_C_R_Z_R,`AO1ANHSX4_C_F_Z_F);
      (B +=> Z) = (`AO1ANHSX4_B_R_Z_R,`AO1ANHSX4_B_F_Z_F);
      (A -=> Z) = (`AO1ANHSX4_A_F_Z_R,`AO1ANHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO1ANHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:39 and Version :1.1 //
 
//  START 
// CELL AO1ANHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1ANHSX8_D_F_Z_F 0.1
`define AO1ANHSX8_D_R_Z_R 0.1
`define AO1ANHSX8_C_F_Z_F 0.1
`define AO1ANHSX8_C_R_Z_R 0.1
`define AO1ANHSX8_B_F_Z_F 0.1
`define AO1ANHSX8_B_R_Z_R 0.1
`define AO1ANHSX8_A_F_Z_R 0.1
`define AO1ANHSX8_A_R_Z_F 0.1

module AO1ANHSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, AndAXB_, C, D);
   and  u1 (AndAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO1ANHSX8_D_R_Z_R,`AO1ANHSX8_D_F_Z_F);
      (C +=> Z) = (`AO1ANHSX8_C_R_Z_R,`AO1ANHSX8_C_F_Z_F);
      (B +=> Z) = (`AO1ANHSX8_B_R_Z_R,`AO1ANHSX8_B_F_Z_F);
      (A -=> Z) = (`AO1ANHSX8_A_F_Z_R,`AO1ANHSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AO1ANHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:39 and Version :1.1 //
 
//  START 
// CELL F_AO1ANHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO1ANHSX4_D_F_Z_F 0.1
`define F_AO1ANHSX4_D_R_Z_R 0.1
`define F_AO1ANHSX4_C_F_Z_F 0.1
`define F_AO1ANHSX4_C_R_Z_R 0.1
`define F_AO1ANHSX4_B_F_Z_F 0.1
`define F_AO1ANHSX4_B_R_Z_R 0.1
`define F_AO1ANHSX4_A_F_Z_R 0.1
`define F_AO1ANHSX4_A_R_Z_F 0.1

module F_AO1ANHSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, AndAXB_, C, D);
   and  u1 (AndAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (D +=> Z) = (`F_AO1ANHSX4_D_R_Z_R,`F_AO1ANHSX4_D_F_Z_F);
      (C +=> Z) = (`F_AO1ANHSX4_C_R_Z_R,`F_AO1ANHSX4_C_F_Z_F);
      (B +=> Z) = (`F_AO1ANHSX4_B_R_Z_R,`F_AO1ANHSX4_B_F_Z_F);
      (A -=> Z) = (`F_AO1ANHSX4_A_F_Z_R,`F_AO1ANHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // F_AO1ANHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:39 and Version :1.1 //
 
//  START 
// CELL AO1CHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1CHS_D_F_Z_R 0.1
`define AO1CHS_D_R_Z_F 0.1
`define AO1CHS_C_F_Z_F 0.1
`define AO1CHS_C_R_Z_R 0.1
`define AO1CHS_B_F_Z_R 0.1
`define AO1CHS_B_R_Z_F 0.1
`define AO1CHS_A_F_Z_R 0.1
`define AO1CHS_A_R_Z_F 0.1

module AO1CHS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAB_, CX, D);
   not  u1 (CX, C);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO1CHS_D_F_Z_R,`AO1CHS_D_R_Z_F);
      (C +=> Z) = (`AO1CHS_C_R_Z_R,`AO1CHS_C_F_Z_F);
      (B -=> Z) = (`AO1CHS_B_F_Z_R,`AO1CHS_B_R_Z_F);
      (A -=> Z) = (`AO1CHS_A_F_Z_R,`AO1CHS_A_R_Z_F);

   endspecify
`endif


endmodule // AO1CHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:46 and Version :1.1 //
 
//  START 
// CELL AO1CHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1CHSP_D_F_Z_R 0.1
`define AO1CHSP_D_R_Z_F 0.1
`define AO1CHSP_C_F_Z_F 0.1
`define AO1CHSP_C_R_Z_R 0.1
`define AO1CHSP_B_F_Z_R 0.1
`define AO1CHSP_B_R_Z_F 0.1
`define AO1CHSP_A_F_Z_R 0.1
`define AO1CHSP_A_R_Z_F 0.1

module AO1CHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAB_, CX, D);
   not  u1 (CX, C);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO1CHSP_D_F_Z_R,`AO1CHSP_D_R_Z_F);
      (C +=> Z) = (`AO1CHSP_C_R_Z_R,`AO1CHSP_C_F_Z_F);
      (B -=> Z) = (`AO1CHSP_B_F_Z_R,`AO1CHSP_B_R_Z_F);
      (A -=> Z) = (`AO1CHSP_A_F_Z_R,`AO1CHSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO1CHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:46 and Version :1.1 //
 
//  START 
// CELL AO1CHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1CHSX4_D_F_Z_R 0.1
`define AO1CHSX4_D_R_Z_F 0.1
`define AO1CHSX4_C_F_Z_F 0.1
`define AO1CHSX4_C_R_Z_R 0.1
`define AO1CHSX4_B_F_Z_R 0.1
`define AO1CHSX4_B_R_Z_F 0.1
`define AO1CHSX4_A_F_Z_R 0.1
`define AO1CHSX4_A_R_Z_F 0.1

module AO1CHSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAB_, CX, D);
   not  u1 (CX, C);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO1CHSX4_D_F_Z_R,`AO1CHSX4_D_R_Z_F);
      (C +=> Z) = (`AO1CHSX4_C_R_Z_R,`AO1CHSX4_C_F_Z_F);
      (B -=> Z) = (`AO1CHSX4_B_F_Z_R,`AO1CHSX4_B_R_Z_F);
      (A -=> Z) = (`AO1CHSX4_A_F_Z_R,`AO1CHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO1CHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:46 and Version :1.1 //
 
//  START 
// CELL AO1CHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1CHSX8_D_F_Z_R 0.1
`define AO1CHSX8_D_R_Z_F 0.1
`define AO1CHSX8_C_F_Z_F 0.1
`define AO1CHSX8_C_R_Z_R 0.1
`define AO1CHSX8_B_F_Z_R 0.1
`define AO1CHSX8_B_R_Z_F 0.1
`define AO1CHSX8_A_F_Z_R 0.1
`define AO1CHSX8_A_R_Z_F 0.1

module AO1CHSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAB_, CX, D);
   not  u1 (CX, C);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO1CHSX8_D_F_Z_R,`AO1CHSX8_D_R_Z_F);
      (C +=> Z) = (`AO1CHSX8_C_R_Z_R,`AO1CHSX8_C_F_Z_F);
      (B -=> Z) = (`AO1CHSX8_B_F_Z_R,`AO1CHSX8_B_R_Z_F);
      (A -=> Z) = (`AO1CHSX8_A_F_Z_R,`AO1CHSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AO1CHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:46 and Version :1.1 //
 
//  START 
// CELL AO1CNHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1CNHS_D_F_Z_F 0.1
`define AO1CNHS_D_R_Z_R 0.1
`define AO1CNHS_C_F_Z_R 0.1
`define AO1CNHS_C_R_Z_F 0.1
`define AO1CNHS_B_F_Z_F 0.1
`define AO1CNHS_B_R_Z_R 0.1
`define AO1CNHS_A_F_Z_F 0.1
`define AO1CNHS_A_R_Z_R 0.1

module AO1CNHS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, AndAB_, CX, D);
   not  u1 (CX, C);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO1CNHS_D_R_Z_R,`AO1CNHS_D_F_Z_F);
      (C -=> Z) = (`AO1CNHS_C_F_Z_R,`AO1CNHS_C_R_Z_F);
      (B +=> Z) = (`AO1CNHS_B_R_Z_R,`AO1CNHS_B_F_Z_F);
      (A +=> Z) = (`AO1CNHS_A_R_Z_R,`AO1CNHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO1CNHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:46 and Version :1.1 //
 
//  START 
// CELL AO1CNHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1CNHSP_D_F_Z_F 0.1
`define AO1CNHSP_D_R_Z_R 0.1
`define AO1CNHSP_C_F_Z_R 0.1
`define AO1CNHSP_C_R_Z_F 0.1
`define AO1CNHSP_B_F_Z_F 0.1
`define AO1CNHSP_B_R_Z_R 0.1
`define AO1CNHSP_A_F_Z_F 0.1
`define AO1CNHSP_A_R_Z_R 0.1

module AO1CNHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, AndAB_, CX, D);
   not  u1 (CX, C);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO1CNHSP_D_R_Z_R,`AO1CNHSP_D_F_Z_F);
      (C -=> Z) = (`AO1CNHSP_C_F_Z_R,`AO1CNHSP_C_R_Z_F);
      (B +=> Z) = (`AO1CNHSP_B_R_Z_R,`AO1CNHSP_B_F_Z_F);
      (A +=> Z) = (`AO1CNHSP_A_R_Z_R,`AO1CNHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO1CNHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:46 and Version :1.1 //
 
//  START 
// CELL AO1CNHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1CNHSX4_D_F_Z_F 0.1
`define AO1CNHSX4_D_R_Z_R 0.1
`define AO1CNHSX4_C_F_Z_R 0.1
`define AO1CNHSX4_C_R_Z_F 0.1
`define AO1CNHSX4_B_F_Z_F 0.1
`define AO1CNHSX4_B_R_Z_R 0.1
`define AO1CNHSX4_A_F_Z_F 0.1
`define AO1CNHSX4_A_R_Z_R 0.1

module AO1CNHSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, AndAB_, CX, D);
   not  u1 (CX, C);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO1CNHSX4_D_R_Z_R,`AO1CNHSX4_D_F_Z_F);
      (C -=> Z) = (`AO1CNHSX4_C_F_Z_R,`AO1CNHSX4_C_R_Z_F);
      (B +=> Z) = (`AO1CNHSX4_B_R_Z_R,`AO1CNHSX4_B_F_Z_F);
      (A +=> Z) = (`AO1CNHSX4_A_R_Z_R,`AO1CNHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO1CNHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:46 and Version :1.1 //
 
//  START 
// CELL AO1CNHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1CNHSX8_D_F_Z_F 0.1
`define AO1CNHSX8_D_R_Z_R 0.1
`define AO1CNHSX8_C_F_Z_R 0.1
`define AO1CNHSX8_C_R_Z_F 0.1
`define AO1CNHSX8_B_F_Z_F 0.1
`define AO1CNHSX8_B_R_Z_R 0.1
`define AO1CNHSX8_A_F_Z_F 0.1
`define AO1CNHSX8_A_R_Z_R 0.1

module AO1CNHSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, AndAB_, CX, D);
   not  u1 (CX, C);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO1CNHSX8_D_R_Z_R,`AO1CNHSX8_D_F_Z_F);
      (C -=> Z) = (`AO1CNHSX8_C_F_Z_R,`AO1CNHSX8_C_R_Z_F);
      (B +=> Z) = (`AO1CNHSX8_B_R_Z_R,`AO1CNHSX8_B_F_Z_F);
      (A +=> Z) = (`AO1CNHSX8_A_R_Z_R,`AO1CNHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO1CNHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:46 and Version :1.1 //
 
//  START 
// CELL AO1NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1NHS_D_F_Z_F 0.1
`define AO1NHS_D_R_Z_R 0.1
`define AO1NHS_C_F_Z_F 0.1
`define AO1NHS_C_R_Z_R 0.1
`define AO1NHS_B_F_Z_F 0.1
`define AO1NHS_B_R_Z_R 0.1
`define AO1NHS_A_F_Z_F 0.1
`define AO1NHS_A_R_Z_R 0.1

module AO1NHS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, AndAB_, C, D);
   and  u1 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO1NHS_D_R_Z_R,`AO1NHS_D_F_Z_F);
      (C +=> Z) = (`AO1NHS_C_R_Z_R,`AO1NHS_C_F_Z_F);
      (B +=> Z) = (`AO1NHS_B_R_Z_R,`AO1NHS_B_F_Z_F);
      (A +=> Z) = (`AO1NHS_A_R_Z_R,`AO1NHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO1NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:49 and Version :1.1 //
 
//  START 
// CELL AO1NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1NHSP_D_F_Z_F 0.1
`define AO1NHSP_D_R_Z_R 0.1
`define AO1NHSP_C_F_Z_F 0.1
`define AO1NHSP_C_R_Z_R 0.1
`define AO1NHSP_B_F_Z_F 0.1
`define AO1NHSP_B_R_Z_R 0.1
`define AO1NHSP_A_F_Z_F 0.1
`define AO1NHSP_A_R_Z_R 0.1

module AO1NHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, AndAB_, C, D);
   and  u1 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO1NHSP_D_R_Z_R,`AO1NHSP_D_F_Z_F);
      (C +=> Z) = (`AO1NHSP_C_R_Z_R,`AO1NHSP_C_F_Z_F);
      (B +=> Z) = (`AO1NHSP_B_R_Z_R,`AO1NHSP_B_F_Z_F);
      (A +=> Z) = (`AO1NHSP_A_R_Z_R,`AO1NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO1NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:49 and Version :1.1 //
 
//  START 
// CELL AO1NHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1NHSX4_D_F_Z_F 0.1
`define AO1NHSX4_D_R_Z_R 0.1
`define AO1NHSX4_C_F_Z_F 0.1
`define AO1NHSX4_C_R_Z_R 0.1
`define AO1NHSX4_B_F_Z_F 0.1
`define AO1NHSX4_B_R_Z_R 0.1
`define AO1NHSX4_A_F_Z_F 0.1
`define AO1NHSX4_A_R_Z_R 0.1

module AO1NHSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, AndAB_, C, D);
   and  u1 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO1NHSX4_D_R_Z_R,`AO1NHSX4_D_F_Z_F);
      (C +=> Z) = (`AO1NHSX4_C_R_Z_R,`AO1NHSX4_C_F_Z_F);
      (B +=> Z) = (`AO1NHSX4_B_R_Z_R,`AO1NHSX4_B_F_Z_F);
      (A +=> Z) = (`AO1NHSX4_A_R_Z_R,`AO1NHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO1NHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:49 and Version :1.1 //
 
//  START 
// CELL AO1NHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO1NHSX8_D_F_Z_F 0.1
`define AO1NHSX8_D_R_Z_R 0.1
`define AO1NHSX8_C_F_Z_F 0.1
`define AO1NHSX8_C_R_Z_R 0.1
`define AO1NHSX8_B_F_Z_F 0.1
`define AO1NHSX8_B_R_Z_R 0.1
`define AO1NHSX8_A_F_Z_F 0.1
`define AO1NHSX8_A_R_Z_R 0.1

module AO1NHSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, AndAB_, C, D);
   and  u1 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO1NHSX8_D_R_Z_R,`AO1NHSX8_D_F_Z_F);
      (C +=> Z) = (`AO1NHSX8_C_R_Z_R,`AO1NHSX8_C_F_Z_F);
      (B +=> Z) = (`AO1NHSX8_B_R_Z_R,`AO1NHSX8_B_F_Z_F);
      (A +=> Z) = (`AO1NHSX8_A_R_Z_R,`AO1NHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO1NHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:49 and Version :1.1 //
 
//  START 
// CELL AO2HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO2HSX05_D_F_Z_R 0.1
`define AO2HSX05_D_R_Z_F 0.1
`define AO2HSX05_C_F_Z_R 0.1
`define AO2HSX05_C_R_Z_F 0.1
`define AO2HSX05_B_F_Z_R 0.1
`define AO2HSX05_B_R_Z_F 0.1
`define AO2HSX05_A_F_Z_R 0.1
`define AO2HSX05_A_R_Z_F 0.1

module AO2HSX05 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAB_, AndCD_);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO2HSX05_D_F_Z_R,`AO2HSX05_D_R_Z_F);
      (C -=> Z) = (`AO2HSX05_C_F_Z_R,`AO2HSX05_C_R_Z_F);
      (B -=> Z) = (`AO2HSX05_B_F_Z_R,`AO2HSX05_B_R_Z_F);
      (A -=> Z) = (`AO2HSX05_A_F_Z_R,`AO2HSX05_A_R_Z_F);

   endspecify
`endif


endmodule  // AO2HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:55 and Version :1.1 //
 
//  START 
// CELL AO2HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO2HS_D_F_Z_R 0.1
`define AO2HS_D_R_Z_F 0.1
`define AO2HS_C_F_Z_R 0.1
`define AO2HS_C_R_Z_F 0.1
`define AO2HS_B_F_Z_R 0.1
`define AO2HS_B_R_Z_F 0.1
`define AO2HS_A_F_Z_R 0.1
`define AO2HS_A_R_Z_F 0.1

module AO2HS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAB_, AndCD_);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO2HS_D_F_Z_R,`AO2HS_D_R_Z_F);
      (C -=> Z) = (`AO2HS_C_F_Z_R,`AO2HS_C_R_Z_F);
      (B -=> Z) = (`AO2HS_B_F_Z_R,`AO2HS_B_R_Z_F);
      (A -=> Z) = (`AO2HS_A_F_Z_R,`AO2HS_A_R_Z_F);

   endspecify
`endif


endmodule  // AO2HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:55 and Version :1.1 //
 
//  START 
// CELL AO2HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO2HSP_D_F_Z_R 0.1
`define AO2HSP_D_R_Z_F 0.1
`define AO2HSP_C_F_Z_R 0.1
`define AO2HSP_C_R_Z_F 0.1
`define AO2HSP_B_F_Z_R 0.1
`define AO2HSP_B_R_Z_F 0.1
`define AO2HSP_A_F_Z_R 0.1
`define AO2HSP_A_R_Z_F 0.1

module AO2HSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAB_, AndCD_);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO2HSP_D_F_Z_R,`AO2HSP_D_R_Z_F);
      (C -=> Z) = (`AO2HSP_C_F_Z_R,`AO2HSP_C_R_Z_F);
      (B -=> Z) = (`AO2HSP_B_F_Z_R,`AO2HSP_B_R_Z_F);
      (A -=> Z) = (`AO2HSP_A_F_Z_R,`AO2HSP_A_R_Z_F);

   endspecify
`endif


endmodule  // AO2HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:55 and Version :1.1 //
 
//  START 
// CELL AO2HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO2HSX4_D_F_Z_R 0.1
`define AO2HSX4_D_R_Z_F 0.1
`define AO2HSX4_C_F_Z_R 0.1
`define AO2HSX4_C_R_Z_F 0.1
`define AO2HSX4_B_F_Z_R 0.1
`define AO2HSX4_B_R_Z_F 0.1
`define AO2HSX4_A_F_Z_R 0.1
`define AO2HSX4_A_R_Z_F 0.1

module AO2HSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAB_, AndCD_);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO2HSX4_D_F_Z_R,`AO2HSX4_D_R_Z_F);
      (C -=> Z) = (`AO2HSX4_C_F_Z_R,`AO2HSX4_C_R_Z_F);
      (B -=> Z) = (`AO2HSX4_B_F_Z_R,`AO2HSX4_B_R_Z_F);
      (A -=> Z) = (`AO2HSX4_A_F_Z_R,`AO2HSX4_A_R_Z_F);

   endspecify
`endif


endmodule  // AO2HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:55 and Version :1.1 //
 
//  START 
// CELL AO2HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO2HSX8_D_F_Z_R 0.1
`define AO2HSX8_D_R_Z_F 0.1
`define AO2HSX8_C_F_Z_R 0.1
`define AO2HSX8_C_R_Z_F 0.1
`define AO2HSX8_B_F_Z_R 0.1
`define AO2HSX8_B_R_Z_F 0.1
`define AO2HSX8_A_F_Z_R 0.1
`define AO2HSX8_A_R_Z_F 0.1

module AO2HSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAB_, AndCD_);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO2HSX8_D_F_Z_R,`AO2HSX8_D_R_Z_F);
      (C -=> Z) = (`AO2HSX8_C_F_Z_R,`AO2HSX8_C_R_Z_F);
      (B -=> Z) = (`AO2HSX8_B_F_Z_R,`AO2HSX8_B_R_Z_F);
      (A -=> Z) = (`AO2HSX8_A_F_Z_R,`AO2HSX8_A_R_Z_F);

   endspecify
`endif


endmodule  // AO2HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:55 and Version :1.1 //
 
//  START 
// CELL F_AO2HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO2HS_D_F_Z_R 0.1
`define F_AO2HS_D_R_Z_F 0.1
`define F_AO2HS_C_F_Z_R 0.1
`define F_AO2HS_C_R_Z_F 0.1
`define F_AO2HS_B_F_Z_R 0.1
`define F_AO2HS_B_R_Z_F 0.1
`define F_AO2HS_A_F_Z_R 0.1
`define F_AO2HS_A_R_Z_F 0.1

module F_AO2HS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAB_, AndCD_);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`F_AO2HS_D_F_Z_R,`F_AO2HS_D_R_Z_F);
      (C -=> Z) = (`F_AO2HS_C_F_Z_R,`F_AO2HS_C_R_Z_F);
      (B -=> Z) = (`F_AO2HS_B_F_Z_R,`F_AO2HS_B_R_Z_F);
      (A -=> Z) = (`F_AO2HS_A_F_Z_R,`F_AO2HS_A_R_Z_F);

   endspecify
`endif


endmodule  // F_AO2HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:55 and Version :1.1 //
 
//  START 
// CELL F_AO2HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO2HSP_D_F_Z_R 0.1
`define F_AO2HSP_D_R_Z_F 0.1
`define F_AO2HSP_C_F_Z_R 0.1
`define F_AO2HSP_C_R_Z_F 0.1
`define F_AO2HSP_B_F_Z_R 0.1
`define F_AO2HSP_B_R_Z_F 0.1
`define F_AO2HSP_A_F_Z_R 0.1
`define F_AO2HSP_A_R_Z_F 0.1

module F_AO2HSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAB_, AndCD_);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`F_AO2HSP_D_F_Z_R,`F_AO2HSP_D_R_Z_F);
      (C -=> Z) = (`F_AO2HSP_C_F_Z_R,`F_AO2HSP_C_R_Z_F);
      (B -=> Z) = (`F_AO2HSP_B_F_Z_R,`F_AO2HSP_B_R_Z_F);
      (A -=> Z) = (`F_AO2HSP_A_F_Z_R,`F_AO2HSP_A_R_Z_F);

   endspecify
`endif


endmodule  // F_AO2HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:05:55 and Version :1.1 //
 
//  START 
// CELL AO20HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO20HSX05_D_F_Z_R 0.1
`define AO20HSX05_D_R_Z_F 0.1
`define AO20HSX05_C_F_Z_R 0.1
`define AO20HSX05_C_R_Z_F 0.1
`define AO20HSX05_B_F_Z_R 0.1
`define AO20HSX05_B_R_Z_F 0.1
`define AO20HSX05_A_F_Z_R 0.1
`define AO20HSX05_A_R_Z_F 0.1

module AO20HSX05 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndOrAB_C_, D);
   and  u1 (AndOrAB_C_, OrAB_, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO20HSX05_D_F_Z_R,`AO20HSX05_D_R_Z_F);
      (C -=> Z) = (`AO20HSX05_C_F_Z_R,`AO20HSX05_C_R_Z_F);
      (B -=> Z) = (`AO20HSX05_B_F_Z_R,`AO20HSX05_B_R_Z_F);
      (A -=> Z) = (`AO20HSX05_A_F_Z_R,`AO20HSX05_A_R_Z_F);

   endspecify
`endif


endmodule  // AO20HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:06:18 and Version :1.1 //
 
//  START 
// CELL AO20HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO20HS_D_F_Z_R 0.1
`define AO20HS_D_R_Z_F 0.1
`define AO20HS_C_F_Z_R 0.1
`define AO20HS_C_R_Z_F 0.1
`define AO20HS_B_F_Z_R 0.1
`define AO20HS_B_R_Z_F 0.1
`define AO20HS_A_F_Z_R 0.1
`define AO20HS_A_R_Z_F 0.1

module AO20HS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndOrAB_C_, D);
   and  u1 (AndOrAB_C_, OrAB_, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO20HS_D_F_Z_R,`AO20HS_D_R_Z_F);
      (C -=> Z) = (`AO20HS_C_F_Z_R,`AO20HS_C_R_Z_F);
      (B -=> Z) = (`AO20HS_B_F_Z_R,`AO20HS_B_R_Z_F);
      (A -=> Z) = (`AO20HS_A_F_Z_R,`AO20HS_A_R_Z_F);

   endspecify
`endif


endmodule  // AO20HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:06:18 and Version :1.1 //
 
//  START 
// CELL AO20HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO20HSP_D_F_Z_R 0.1
`define AO20HSP_D_R_Z_F 0.1
`define AO20HSP_C_F_Z_R 0.1
`define AO20HSP_C_R_Z_F 0.1
`define AO20HSP_B_F_Z_R 0.1
`define AO20HSP_B_R_Z_F 0.1
`define AO20HSP_A_F_Z_R 0.1
`define AO20HSP_A_R_Z_F 0.1

module AO20HSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndOrAB_C_, D);
   and  u1 (AndOrAB_C_, OrAB_, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO20HSP_D_F_Z_R,`AO20HSP_D_R_Z_F);
      (C -=> Z) = (`AO20HSP_C_F_Z_R,`AO20HSP_C_R_Z_F);
      (B -=> Z) = (`AO20HSP_B_F_Z_R,`AO20HSP_B_R_Z_F);
      (A -=> Z) = (`AO20HSP_A_F_Z_R,`AO20HSP_A_R_Z_F);

   endspecify
`endif


endmodule  // AO20HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:06:18 and Version :1.1 //
 
//  START 
// CELL AO20HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO20HSX4_D_F_Z_R 0.1
`define AO20HSX4_D_R_Z_F 0.1
`define AO20HSX4_C_F_Z_R 0.1
`define AO20HSX4_C_R_Z_F 0.1
`define AO20HSX4_B_F_Z_R 0.1
`define AO20HSX4_B_R_Z_F 0.1
`define AO20HSX4_A_F_Z_R 0.1
`define AO20HSX4_A_R_Z_F 0.1

module AO20HSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndOrAB_C_, D);
   and  u1 (AndOrAB_C_, OrAB_, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO20HSX4_D_F_Z_R,`AO20HSX4_D_R_Z_F);
      (C -=> Z) = (`AO20HSX4_C_F_Z_R,`AO20HSX4_C_R_Z_F);
      (B -=> Z) = (`AO20HSX4_B_F_Z_R,`AO20HSX4_B_R_Z_F);
      (A -=> Z) = (`AO20HSX4_A_F_Z_R,`AO20HSX4_A_R_Z_F);

   endspecify
`endif


endmodule  // AO20HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:06:18 and Version :1.1 //
 
//  START 
// CELL AO20HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO20HSX8_D_F_Z_R 0.1
`define AO20HSX8_D_R_Z_F 0.1
`define AO20HSX8_C_F_Z_R 0.1
`define AO20HSX8_C_R_Z_F 0.1
`define AO20HSX8_B_F_Z_R 0.1
`define AO20HSX8_B_R_Z_F 0.1
`define AO20HSX8_A_F_Z_R 0.1
`define AO20HSX8_A_R_Z_F 0.1

module AO20HSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndOrAB_C_, D);
   and  u1 (AndOrAB_C_, OrAB_, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO20HSX8_D_F_Z_R,`AO20HSX8_D_R_Z_F);
      (C -=> Z) = (`AO20HSX8_C_F_Z_R,`AO20HSX8_C_R_Z_F);
      (B -=> Z) = (`AO20HSX8_B_F_Z_R,`AO20HSX8_B_R_Z_F);
      (A -=> Z) = (`AO20HSX8_A_F_Z_R,`AO20HSX8_A_R_Z_F);

   endspecify
`endif


endmodule  // AO20HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:06:18 and Version :1.1 //
 
//  START 
// CELL AO20NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO20NHS_D_F_Z_F 0.1
`define AO20NHS_D_R_Z_R 0.1
`define AO20NHS_C_F_Z_F 0.1
`define AO20NHS_C_R_Z_R 0.1
`define AO20NHS_B_F_Z_F 0.1
`define AO20NHS_B_R_Z_R 0.1
`define AO20NHS_A_F_Z_F 0.1
`define AO20NHS_A_R_Z_R 0.1

module AO20NHS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (OrAB_, A, B);
   and  u1 (AndOrAB_C_, OrAB_, C);
   or  u2 (Z, AndOrAB_C_, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO20NHS_D_R_Z_R,`AO20NHS_D_F_Z_F);
      (C +=> Z) = (`AO20NHS_C_R_Z_R,`AO20NHS_C_F_Z_F);
      (B +=> Z) = (`AO20NHS_B_R_Z_R,`AO20NHS_B_F_Z_F);
      (A +=> Z) = (`AO20NHS_A_R_Z_R,`AO20NHS_A_F_Z_F);

   endspecify
`endif


endmodule  // AO20NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:06:18 and Version :1.1 //
 
//  START 
// CELL AO20NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO20NHSP_D_F_Z_F 0.1
`define AO20NHSP_D_R_Z_R 0.1
`define AO20NHSP_C_F_Z_F 0.1
`define AO20NHSP_C_R_Z_R 0.1
`define AO20NHSP_B_F_Z_F 0.1
`define AO20NHSP_B_R_Z_R 0.1
`define AO20NHSP_A_F_Z_F 0.1
`define AO20NHSP_A_R_Z_R 0.1

module AO20NHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (OrAB_, A, B);
   and  u1 (AndOrAB_C_, OrAB_, C);
   or  u2 (Z, AndOrAB_C_, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO20NHSP_D_R_Z_R,`AO20NHSP_D_F_Z_F);
      (C +=> Z) = (`AO20NHSP_C_R_Z_R,`AO20NHSP_C_F_Z_F);
      (B +=> Z) = (`AO20NHSP_B_R_Z_R,`AO20NHSP_B_F_Z_F);
      (A +=> Z) = (`AO20NHSP_A_R_Z_R,`AO20NHSP_A_F_Z_F);

   endspecify
`endif


endmodule  // AO20NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:06:18 and Version :1.1 //
 
//  START 
// CELL AO20NHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO20NHSX4_D_F_Z_F 0.1
`define AO20NHSX4_D_R_Z_R 0.1
`define AO20NHSX4_C_F_Z_F 0.1
`define AO20NHSX4_C_R_Z_R 0.1
`define AO20NHSX4_B_F_Z_F 0.1
`define AO20NHSX4_B_R_Z_R 0.1
`define AO20NHSX4_A_F_Z_F 0.1
`define AO20NHSX4_A_R_Z_R 0.1

module AO20NHSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (OrAB_, A, B);
   and  u1 (AndOrAB_C_, OrAB_, C);
   or  u2 (Z, AndOrAB_C_, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO20NHSX4_D_R_Z_R,`AO20NHSX4_D_F_Z_F);
      (C +=> Z) = (`AO20NHSX4_C_R_Z_R,`AO20NHSX4_C_F_Z_F);
      (B +=> Z) = (`AO20NHSX4_B_R_Z_R,`AO20NHSX4_B_F_Z_F);
      (A +=> Z) = (`AO20NHSX4_A_R_Z_R,`AO20NHSX4_A_F_Z_F);

   endspecify
`endif


endmodule  // AO20NHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:06:18 and Version :1.1 //
 
//  START 
// CELL AO20NHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO20NHSX8_D_F_Z_F 0.1
`define AO20NHSX8_D_R_Z_R 0.1
`define AO20NHSX8_C_F_Z_F 0.1
`define AO20NHSX8_C_R_Z_R 0.1
`define AO20NHSX8_B_F_Z_F 0.1
`define AO20NHSX8_B_R_Z_R 0.1
`define AO20NHSX8_A_F_Z_F 0.1
`define AO20NHSX8_A_R_Z_R 0.1

module AO20NHSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (OrAB_, A, B);
   and  u1 (AndOrAB_C_, OrAB_, C);
   or  u2 (Z, AndOrAB_C_, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO20NHSX8_D_R_Z_R,`AO20NHSX8_D_F_Z_F);
      (C +=> Z) = (`AO20NHSX8_C_R_Z_R,`AO20NHSX8_C_F_Z_F);
      (B +=> Z) = (`AO20NHSX8_B_R_Z_R,`AO20NHSX8_B_F_Z_F);
      (A +=> Z) = (`AO20NHSX8_A_R_Z_R,`AO20NHSX8_A_F_Z_F);

   endspecify
`endif


endmodule  // AO20NHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:06:18 and Version :1.1 //
 
//  START 
// CELL AO21HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO21HSX05_D_F_Z_R 0.1
`define AO21HSX05_D_R_Z_F 0.1
`define AO21HSX05_C_F_Z_R 0.1
`define AO21HSX05_C_R_Z_F 0.1
`define AO21HSX05_B_F_Z_R 0.1
`define AO21HSX05_B_R_Z_F 0.1
`define AO21HSX05_A_F_Z_R 0.1
`define AO21HSX05_A_R_Z_F 0.1

module AO21HSX05 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrABC_, D);
   or  u1 (OrABC_, A, B, C);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO21HSX05_D_F_Z_R,`AO21HSX05_D_R_Z_F);
      (C -=> Z) = (`AO21HSX05_C_F_Z_R,`AO21HSX05_C_R_Z_F);
      (B -=> Z) = (`AO21HSX05_B_F_Z_R,`AO21HSX05_B_R_Z_F);
      (A -=> Z) = (`AO21HSX05_A_F_Z_R,`AO21HSX05_A_R_Z_F);

   endspecify
`endif


endmodule  // AO21HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:06:37 and Version :1.1 //
 
//  START 
// CELL AO21HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO21HS_D_F_Z_R 0.1
`define AO21HS_D_R_Z_F 0.1
`define AO21HS_C_F_Z_R 0.1
`define AO21HS_C_R_Z_F 0.1
`define AO21HS_B_F_Z_R 0.1
`define AO21HS_B_R_Z_F 0.1
`define AO21HS_A_F_Z_R 0.1
`define AO21HS_A_R_Z_F 0.1

module AO21HS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrABC_, D);
   or  u1 (OrABC_, A, B, C);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO21HS_D_F_Z_R,`AO21HS_D_R_Z_F);
      (C -=> Z) = (`AO21HS_C_F_Z_R,`AO21HS_C_R_Z_F);
      (B -=> Z) = (`AO21HS_B_F_Z_R,`AO21HS_B_R_Z_F);
      (A -=> Z) = (`AO21HS_A_F_Z_R,`AO21HS_A_R_Z_F);

   endspecify
`endif


endmodule  // AO21HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:06:37 and Version :1.1 //
 
//  START 
// CELL AO21HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO21HSP_D_F_Z_R 0.1
`define AO21HSP_D_R_Z_F 0.1
`define AO21HSP_C_F_Z_R 0.1
`define AO21HSP_C_R_Z_F 0.1
`define AO21HSP_B_F_Z_R 0.1
`define AO21HSP_B_R_Z_F 0.1
`define AO21HSP_A_F_Z_R 0.1
`define AO21HSP_A_R_Z_F 0.1

module AO21HSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrABC_, D);
   or  u1 (OrABC_, A, B, C);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO21HSP_D_F_Z_R,`AO21HSP_D_R_Z_F);
      (C -=> Z) = (`AO21HSP_C_F_Z_R,`AO21HSP_C_R_Z_F);
      (B -=> Z) = (`AO21HSP_B_F_Z_R,`AO21HSP_B_R_Z_F);
      (A -=> Z) = (`AO21HSP_A_F_Z_R,`AO21HSP_A_R_Z_F);

   endspecify
`endif


endmodule  // AO21HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:06:37 and Version :1.1 //
 
//  START 
// CELL AO21NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO21NHS_D_F_Z_F 0.1
`define AO21NHS_D_R_Z_R 0.1
`define AO21NHS_C_F_Z_F 0.1
`define AO21NHS_C_R_Z_R 0.1
`define AO21NHS_B_F_Z_F 0.1
`define AO21NHS_B_R_Z_R 0.1
`define AO21NHS_A_F_Z_F 0.1
`define AO21NHS_A_R_Z_R 0.1

module AO21NHS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (OrABC_, A, B, C);
   and  u1 (Z, OrABC_, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO21NHS_D_R_Z_R,`AO21NHS_D_F_Z_F);
      (C +=> Z) = (`AO21NHS_C_R_Z_R,`AO21NHS_C_F_Z_F);
      (B +=> Z) = (`AO21NHS_B_R_Z_R,`AO21NHS_B_F_Z_F);
      (A +=> Z) = (`AO21NHS_A_R_Z_R,`AO21NHS_A_F_Z_F);

   endspecify
`endif


endmodule  // AO21NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:06:37 and Version :1.1 //
 
//  START 
// CELL AO21NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO21NHSP_D_F_Z_F 0.1
`define AO21NHSP_D_R_Z_R 0.1
`define AO21NHSP_C_F_Z_F 0.1
`define AO21NHSP_C_R_Z_R 0.1
`define AO21NHSP_B_F_Z_F 0.1
`define AO21NHSP_B_R_Z_R 0.1
`define AO21NHSP_A_F_Z_F 0.1
`define AO21NHSP_A_R_Z_R 0.1

module AO21NHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (OrABC_, A, B, C);
   and  u1 (Z, OrABC_, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO21NHSP_D_R_Z_R,`AO21NHSP_D_F_Z_F);
      (C +=> Z) = (`AO21NHSP_C_R_Z_R,`AO21NHSP_C_F_Z_F);
      (B +=> Z) = (`AO21NHSP_B_R_Z_R,`AO21NHSP_B_F_Z_F);
      (A +=> Z) = (`AO21NHSP_A_R_Z_R,`AO21NHSP_A_F_Z_F);

   endspecify
`endif


endmodule  // AO21NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:06:37 and Version :1.1 //
 
//  START 
// CELL AO21NHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO21NHSX4_D_F_Z_F 0.1
`define AO21NHSX4_D_R_Z_R 0.1
`define AO21NHSX4_C_F_Z_F 0.1
`define AO21NHSX4_C_R_Z_R 0.1
`define AO21NHSX4_B_F_Z_F 0.1
`define AO21NHSX4_B_R_Z_R 0.1
`define AO21NHSX4_A_F_Z_F 0.1
`define AO21NHSX4_A_R_Z_R 0.1

module AO21NHSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (OrABC_, A, B, C);
   and  u1 (Z, OrABC_, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO21NHSX4_D_R_Z_R,`AO21NHSX4_D_F_Z_F);
      (C +=> Z) = (`AO21NHSX4_C_R_Z_R,`AO21NHSX4_C_F_Z_F);
      (B +=> Z) = (`AO21NHSX4_B_R_Z_R,`AO21NHSX4_B_F_Z_F);
      (A +=> Z) = (`AO21NHSX4_A_R_Z_R,`AO21NHSX4_A_F_Z_F);

   endspecify
`endif


endmodule  // AO21NHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:06:37 and Version :1.1 //
 
//  START 
// CELL AO22HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO22HSX05_E_F_Z_R 0.1
`define AO22HSX05_E_R_Z_F 0.1
`define AO22HSX05_D_F_Z_R 0.1
`define AO22HSX05_D_R_Z_F 0.1
`define AO22HSX05_C_F_Z_R 0.1
`define AO22HSX05_C_R_Z_F 0.1
`define AO22HSX05_B_F_Z_R 0.1
`define AO22HSX05_B_R_Z_F 0.1
`define AO22HSX05_A_F_Z_R 0.1
`define AO22HSX05_A_R_Z_F 0.1

module AO22HSX05 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   nand  u0 (Z, OrABC_, OrDE_);
   or  u1 (OrDE_, D, E);
   or  u2 (OrABC_, A, B, C);


`ifdef functional
`else
   specify

      (E -=> Z) = (`AO22HSX05_E_F_Z_R,`AO22HSX05_E_R_Z_F);
      (D -=> Z) = (`AO22HSX05_D_F_Z_R,`AO22HSX05_D_R_Z_F);
      (C -=> Z) = (`AO22HSX05_C_F_Z_R,`AO22HSX05_C_R_Z_F);
      (B -=> Z) = (`AO22HSX05_B_F_Z_R,`AO22HSX05_B_R_Z_F);
      (A -=> Z) = (`AO22HSX05_A_F_Z_R,`AO22HSX05_A_R_Z_F);

   endspecify
`endif


endmodule  // AO22HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:06:56 and Version :1.1 //
 
//  START 
// CELL AO22HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO22HS_E_F_Z_R 0.1
`define AO22HS_E_R_Z_F 0.1
`define AO22HS_D_F_Z_R 0.1
`define AO22HS_D_R_Z_F 0.1
`define AO22HS_C_F_Z_R 0.1
`define AO22HS_C_R_Z_F 0.1
`define AO22HS_B_F_Z_R 0.1
`define AO22HS_B_R_Z_F 0.1
`define AO22HS_A_F_Z_R 0.1
`define AO22HS_A_R_Z_F 0.1

module AO22HS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   nand  u0 (Z, OrABC_, OrDE_);
   or  u1 (OrDE_, D, E);
   or  u2 (OrABC_, A, B, C);


`ifdef functional
`else
   specify

      (E -=> Z) = (`AO22HS_E_F_Z_R,`AO22HS_E_R_Z_F);
      (D -=> Z) = (`AO22HS_D_F_Z_R,`AO22HS_D_R_Z_F);
      (C -=> Z) = (`AO22HS_C_F_Z_R,`AO22HS_C_R_Z_F);
      (B -=> Z) = (`AO22HS_B_F_Z_R,`AO22HS_B_R_Z_F);
      (A -=> Z) = (`AO22HS_A_F_Z_R,`AO22HS_A_R_Z_F);

   endspecify
`endif


endmodule  // AO22HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:06:56 and Version :1.1 //
 
//  START 
// CELL AO22NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO22NHS_E_F_Z_F 0.1
`define AO22NHS_E_R_Z_R 0.1
`define AO22NHS_D_F_Z_F 0.1
`define AO22NHS_D_R_Z_R 0.1
`define AO22NHS_C_F_Z_F 0.1
`define AO22NHS_C_R_Z_R 0.1
`define AO22NHS_B_F_Z_F 0.1
`define AO22NHS_B_R_Z_R 0.1
`define AO22NHS_A_F_Z_F 0.1
`define AO22NHS_A_R_Z_R 0.1

module AO22NHS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   or  u0 (OrABC_, A, B, C);
   or  u1 (OrDE_, D, E);
   and  u2 (Z, OrABC_, OrDE_);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO22NHS_E_R_Z_R,`AO22NHS_E_F_Z_F);
      (D +=> Z) = (`AO22NHS_D_R_Z_R,`AO22NHS_D_F_Z_F);
      (C +=> Z) = (`AO22NHS_C_R_Z_R,`AO22NHS_C_F_Z_F);
      (B +=> Z) = (`AO22NHS_B_R_Z_R,`AO22NHS_B_F_Z_F);
      (A +=> Z) = (`AO22NHS_A_R_Z_R,`AO22NHS_A_F_Z_F);

   endspecify
`endif


endmodule  // AO22NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:06:56 and Version :1.1 //
 
//  START 
// CELL AO22NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO22NHSP_E_F_Z_F 0.1
`define AO22NHSP_E_R_Z_R 0.1
`define AO22NHSP_D_F_Z_F 0.1
`define AO22NHSP_D_R_Z_R 0.1
`define AO22NHSP_C_F_Z_F 0.1
`define AO22NHSP_C_R_Z_R 0.1
`define AO22NHSP_B_F_Z_F 0.1
`define AO22NHSP_B_R_Z_R 0.1
`define AO22NHSP_A_F_Z_F 0.1
`define AO22NHSP_A_R_Z_R 0.1

module AO22NHSP (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   or  u0 (OrABC_, A, B, C);
   or  u1 (OrDE_, D, E);
   and  u2 (Z, OrABC_, OrDE_);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO22NHSP_E_R_Z_R,`AO22NHSP_E_F_Z_F);
      (D +=> Z) = (`AO22NHSP_D_R_Z_R,`AO22NHSP_D_F_Z_F);
      (C +=> Z) = (`AO22NHSP_C_R_Z_R,`AO22NHSP_C_F_Z_F);
      (B +=> Z) = (`AO22NHSP_B_R_Z_R,`AO22NHSP_B_F_Z_F);
      (A +=> Z) = (`AO22NHSP_A_R_Z_R,`AO22NHSP_A_F_Z_F);

   endspecify
`endif


endmodule  // AO22NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:06:56 and Version :1.1 //
 
//  START 
// CELL AO23HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO23HSX05_E_F_Z_R 0.1
`define AO23HSX05_E_R_Z_F 0.1
`define AO23HSX05_D_F_Z_R 0.1
`define AO23HSX05_D_R_Z_F 0.1
`define AO23HSX05_C_F_Z_R 0.1
`define AO23HSX05_C_R_Z_F 0.1
`define AO23HSX05_B_F_Z_R 0.1
`define AO23HSX05_B_R_Z_F 0.1
`define AO23HSX05_A_F_Z_R 0.1
`define AO23HSX05_A_R_Z_F 0.1

module AO23HSX05 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   or  u0 (OrAB_, A, B);
   or  u1 (OrCD_, C, D);
   nand  u2 (Z, OrAB_, OrCD_, E);


`ifdef functional
`else
   specify

      (E -=> Z) = (`AO23HSX05_E_F_Z_R,`AO23HSX05_E_R_Z_F);
      (D -=> Z) = (`AO23HSX05_D_F_Z_R,`AO23HSX05_D_R_Z_F);
      (C -=> Z) = (`AO23HSX05_C_F_Z_R,`AO23HSX05_C_R_Z_F);
      (B -=> Z) = (`AO23HSX05_B_F_Z_R,`AO23HSX05_B_R_Z_F);
      (A -=> Z) = (`AO23HSX05_A_F_Z_R,`AO23HSX05_A_R_Z_F);

   endspecify
`endif


endmodule  // AO23HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:07:15 and Version :1.1 //
 
//  START 
// CELL AO23HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO23HS_E_F_Z_R 0.1
`define AO23HS_E_R_Z_F 0.1
`define AO23HS_D_F_Z_R 0.1
`define AO23HS_D_R_Z_F 0.1
`define AO23HS_C_F_Z_R 0.1
`define AO23HS_C_R_Z_F 0.1
`define AO23HS_B_F_Z_R 0.1
`define AO23HS_B_R_Z_F 0.1
`define AO23HS_A_F_Z_R 0.1
`define AO23HS_A_R_Z_F 0.1

module AO23HS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   or  u0 (OrAB_, A, B);
   or  u1 (OrCD_, C, D);
   nand  u2 (Z, OrAB_, OrCD_, E);


`ifdef functional
`else
   specify

      (E -=> Z) = (`AO23HS_E_F_Z_R,`AO23HS_E_R_Z_F);
      (D -=> Z) = (`AO23HS_D_F_Z_R,`AO23HS_D_R_Z_F);
      (C -=> Z) = (`AO23HS_C_F_Z_R,`AO23HS_C_R_Z_F);
      (B -=> Z) = (`AO23HS_B_F_Z_R,`AO23HS_B_R_Z_F);
      (A -=> Z) = (`AO23HS_A_F_Z_R,`AO23HS_A_R_Z_F);

   endspecify
`endif


endmodule  // AO23HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:07:15 and Version :1.1 //
 
//  START 
// CELL AO23NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO23NHS_E_F_Z_F 0.1
`define AO23NHS_E_R_Z_R 0.1
`define AO23NHS_D_F_Z_F 0.1
`define AO23NHS_D_R_Z_R 0.1
`define AO23NHS_C_F_Z_F 0.1
`define AO23NHS_C_R_Z_R 0.1
`define AO23NHS_B_F_Z_F 0.1
`define AO23NHS_B_R_Z_R 0.1
`define AO23NHS_A_F_Z_F 0.1
`define AO23NHS_A_R_Z_R 0.1

module AO23NHS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   or  u0 (OrAB_, A, B);
   or  u1 (OrCD_, C, D);
   and  u2 (Z, OrAB_, OrCD_, E);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO23NHS_E_R_Z_R,`AO23NHS_E_F_Z_F);
      (D +=> Z) = (`AO23NHS_D_R_Z_R,`AO23NHS_D_F_Z_F);
      (C +=> Z) = (`AO23NHS_C_R_Z_R,`AO23NHS_C_F_Z_F);
      (B +=> Z) = (`AO23NHS_B_R_Z_R,`AO23NHS_B_F_Z_F);
      (A +=> Z) = (`AO23NHS_A_R_Z_R,`AO23NHS_A_F_Z_F);

   endspecify
`endif


endmodule  // AO23NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:07:15 and Version :1.1 //
 
//  START 
// CELL AO23NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO23NHSP_E_F_Z_F 0.1
`define AO23NHSP_E_R_Z_R 0.1
`define AO23NHSP_D_F_Z_F 0.1
`define AO23NHSP_D_R_Z_R 0.1
`define AO23NHSP_C_F_Z_F 0.1
`define AO23NHSP_C_R_Z_R 0.1
`define AO23NHSP_B_F_Z_F 0.1
`define AO23NHSP_B_R_Z_R 0.1
`define AO23NHSP_A_F_Z_F 0.1
`define AO23NHSP_A_R_Z_R 0.1

module AO23NHSP (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   or  u0 (OrAB_, A, B);
   or  u1 (OrCD_, C, D);
   and  u2 (Z, OrAB_, OrCD_, E);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO23NHSP_E_R_Z_R,`AO23NHSP_E_F_Z_F);
      (D +=> Z) = (`AO23NHSP_D_R_Z_R,`AO23NHSP_D_F_Z_F);
      (C +=> Z) = (`AO23NHSP_C_R_Z_R,`AO23NHSP_C_F_Z_F);
      (B +=> Z) = (`AO23NHSP_B_R_Z_R,`AO23NHSP_B_F_Z_F);
      (A +=> Z) = (`AO23NHSP_A_R_Z_R,`AO23NHSP_A_F_Z_F);

   endspecify
`endif


endmodule  // AO23NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:07:15 and Version :1.1 //
 
//  START 
// CELL AO24HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO24HSX05_E_F_Z_R 0.1
`define AO24HSX05_E_R_Z_F 0.1
`define AO24HSX05_D_F_Z_R 0.1
`define AO24HSX05_D_R_Z_F 0.1
`define AO24HSX05_C_F_Z_R 0.1
`define AO24HSX05_C_R_Z_F 0.1
`define AO24HSX05_B_F_Z_R 0.1
`define AO24HSX05_B_R_Z_F 0.1
`define AO24HSX05_A_F_Z_R 0.1
`define AO24HSX05_A_R_Z_F 0.1

module AO24HSX05 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   nor  u0 (Z, AndABC_, D, E);
   and  u1 (AndABC_, A, B, C);


`ifdef functional
`else
   specify

      (E -=> Z) = (`AO24HSX05_E_F_Z_R,`AO24HSX05_E_R_Z_F);
      (D -=> Z) = (`AO24HSX05_D_F_Z_R,`AO24HSX05_D_R_Z_F);
      (C -=> Z) = (`AO24HSX05_C_F_Z_R,`AO24HSX05_C_R_Z_F);
      (B -=> Z) = (`AO24HSX05_B_F_Z_R,`AO24HSX05_B_R_Z_F);
      (A -=> Z) = (`AO24HSX05_A_F_Z_R,`AO24HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // AO24HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:07:34 and Version :1.1 //
 
//  START 
// CELL AO24HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO24HS_E_F_Z_R 0.1
`define AO24HS_E_R_Z_F 0.1
`define AO24HS_D_F_Z_R 0.1
`define AO24HS_D_R_Z_F 0.1
`define AO24HS_C_F_Z_R 0.1
`define AO24HS_C_R_Z_F 0.1
`define AO24HS_B_F_Z_R 0.1
`define AO24HS_B_R_Z_F 0.1
`define AO24HS_A_F_Z_R 0.1
`define AO24HS_A_R_Z_F 0.1

module AO24HS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   nor  u0 (Z, AndABC_, D, E);
   and  u1 (AndABC_, A, B, C);


`ifdef functional
`else
   specify

      (E -=> Z) = (`AO24HS_E_F_Z_R,`AO24HS_E_R_Z_F);
      (D -=> Z) = (`AO24HS_D_F_Z_R,`AO24HS_D_R_Z_F);
      (C -=> Z) = (`AO24HS_C_F_Z_R,`AO24HS_C_R_Z_F);
      (B -=> Z) = (`AO24HS_B_F_Z_R,`AO24HS_B_R_Z_F);
      (A -=> Z) = (`AO24HS_A_F_Z_R,`AO24HS_A_R_Z_F);

   endspecify
`endif


endmodule // AO24HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:07:34 and Version :1.1 //
 
//  START 
// CELL AO24NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO24NHS_E_F_Z_F 0.1
`define AO24NHS_E_R_Z_R 0.1
`define AO24NHS_D_F_Z_F 0.1
`define AO24NHS_D_R_Z_R 0.1
`define AO24NHS_C_F_Z_F 0.1
`define AO24NHS_C_R_Z_R 0.1
`define AO24NHS_B_F_Z_F 0.1
`define AO24NHS_B_R_Z_R 0.1
`define AO24NHS_A_F_Z_F 0.1
`define AO24NHS_A_R_Z_R 0.1

module AO24NHS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndABC_, A, B, C);
   or  u1 (Z, AndABC_, D, E);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO24NHS_E_R_Z_R,`AO24NHS_E_F_Z_F);
      (D +=> Z) = (`AO24NHS_D_R_Z_R,`AO24NHS_D_F_Z_F);
      (C +=> Z) = (`AO24NHS_C_R_Z_R,`AO24NHS_C_F_Z_F);
      (B +=> Z) = (`AO24NHS_B_R_Z_R,`AO24NHS_B_F_Z_F);
      (A +=> Z) = (`AO24NHS_A_R_Z_R,`AO24NHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO24NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:07:34 and Version :1.1 //
 
//  START 
// CELL AO24NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO24NHSP_E_F_Z_F 0.1
`define AO24NHSP_E_R_Z_R 0.1
`define AO24NHSP_D_F_Z_F 0.1
`define AO24NHSP_D_R_Z_R 0.1
`define AO24NHSP_C_F_Z_F 0.1
`define AO24NHSP_C_R_Z_R 0.1
`define AO24NHSP_B_F_Z_F 0.1
`define AO24NHSP_B_R_Z_R 0.1
`define AO24NHSP_A_F_Z_F 0.1
`define AO24NHSP_A_R_Z_R 0.1

module AO24NHSP (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndABC_, A, B, C);
   or  u1 (Z, AndABC_, D, E);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO24NHSP_E_R_Z_R,`AO24NHSP_E_F_Z_F);
      (D +=> Z) = (`AO24NHSP_D_R_Z_R,`AO24NHSP_D_F_Z_F);
      (C +=> Z) = (`AO24NHSP_C_R_Z_R,`AO24NHSP_C_F_Z_F);
      (B +=> Z) = (`AO24NHSP_B_R_Z_R,`AO24NHSP_B_F_Z_F);
      (A +=> Z) = (`AO24NHSP_A_R_Z_R,`AO24NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO24NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:07:34 and Version :1.1 //
 
//  START 
// CELL AO25HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO25HS_E_F_Z_R 0.1
`define AO25HS_E_R_Z_F 0.1
`define AO25HS_D_F_Z_R 0.1
`define AO25HS_D_R_Z_F 0.1
`define AO25HS_C_F_Z_R 0.1
`define AO25HS_C_R_Z_F 0.1
`define AO25HS_B_F_Z_R 0.1
`define AO25HS_B_R_Z_F 0.1
`define AO25HS_A_F_Z_R 0.1
`define AO25HS_A_R_Z_F 0.1

module AO25HS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndAB_, A, B);
   or  u1 (OrAndAB_C_, AndAB_, C);
   or  u2 (OrDE_, D, E);
   nand  u3 (Z, OrAndAB_C_, OrDE_);


`ifdef functional
`else
   specify

      (E -=> Z) = (`AO25HS_E_F_Z_R,`AO25HS_E_R_Z_F);
      (D -=> Z) = (`AO25HS_D_F_Z_R,`AO25HS_D_R_Z_F);
      (C -=> Z) = (`AO25HS_C_F_Z_R,`AO25HS_C_R_Z_F);
      (B -=> Z) = (`AO25HS_B_F_Z_R,`AO25HS_B_R_Z_F);
      (A -=> Z) = (`AO25HS_A_F_Z_R,`AO25HS_A_R_Z_F);

   endspecify
`endif


endmodule // AO25HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:07:59 and Version :1.1 //
 
//  START 
// CELL AO25NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO25NHS_E_F_Z_F 0.1
`define AO25NHS_E_R_Z_R 0.1
`define AO25NHS_D_F_Z_F 0.1
`define AO25NHS_D_R_Z_R 0.1
`define AO25NHS_C_F_Z_F 0.1
`define AO25NHS_C_R_Z_R 0.1
`define AO25NHS_B_F_Z_F 0.1
`define AO25NHS_B_R_Z_R 0.1
`define AO25NHS_A_F_Z_F 0.1
`define AO25NHS_A_R_Z_R 0.1

module AO25NHS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndAB_, A, B);
   or  u1 (OrAndAB_C_, AndAB_, C);
   or  u2 (OrDE_, D, E);
   and  u3 (Z, OrAndAB_C_, OrDE_);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO25NHS_E_R_Z_R,`AO25NHS_E_F_Z_F);
      (D +=> Z) = (`AO25NHS_D_R_Z_R,`AO25NHS_D_F_Z_F);
      (C +=> Z) = (`AO25NHS_C_R_Z_R,`AO25NHS_C_F_Z_F);
      (B +=> Z) = (`AO25NHS_B_R_Z_R,`AO25NHS_B_F_Z_F);
      (A +=> Z) = (`AO25NHS_A_R_Z_R,`AO25NHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO25NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:07:59 and Version :1.1 //
 
//  START 
// CELL AO25NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO25NHSP_E_F_Z_F 0.1
`define AO25NHSP_E_R_Z_R 0.1
`define AO25NHSP_D_F_Z_F 0.1
`define AO25NHSP_D_R_Z_R 0.1
`define AO25NHSP_C_F_Z_F 0.1
`define AO25NHSP_C_R_Z_R 0.1
`define AO25NHSP_B_F_Z_F 0.1
`define AO25NHSP_B_R_Z_R 0.1
`define AO25NHSP_A_F_Z_F 0.1
`define AO25NHSP_A_R_Z_R 0.1

module AO25NHSP (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndAB_, A, B);
   or  u1 (OrAndAB_C_, AndAB_, C);
   or  u2 (OrDE_, D, E);
   and  u3 (Z, OrAndAB_C_, OrDE_);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO25NHSP_E_R_Z_R,`AO25NHSP_E_F_Z_F);
      (D +=> Z) = (`AO25NHSP_D_R_Z_R,`AO25NHSP_D_F_Z_F);
      (C +=> Z) = (`AO25NHSP_C_R_Z_R,`AO25NHSP_C_F_Z_F);
      (B +=> Z) = (`AO25NHSP_B_R_Z_R,`AO25NHSP_B_F_Z_F);
      (A +=> Z) = (`AO25NHSP_A_R_Z_R,`AO25NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO25NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:07:59 and Version :1.1 //
 
//  START 
// CELL AO26HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO26HSX05_E_F_Z_R 0.1
`define AO26HSX05_E_R_Z_F 0.1
`define AO26HSX05_D_F_Z_R 0.1
`define AO26HSX05_D_R_Z_F 0.1
`define AO26HSX05_C_F_Z_R 0.1
`define AO26HSX05_C_R_Z_F 0.1
`define AO26HSX05_B_F_Z_R 0.1
`define AO26HSX05_B_R_Z_F 0.1
`define AO26HSX05_A_F_Z_R 0.1
`define AO26HSX05_A_R_Z_F 0.1

module AO26HSX05 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndAB_, A, B);
   or  u1 (OrAndAB_CD_, AndAB_, C, D);
   nand  u2 (Z, OrAndAB_CD_, E);


`ifdef functional
`else
   specify

      (E -=> Z) = (`AO26HSX05_E_F_Z_R,`AO26HSX05_E_R_Z_F);
      (D -=> Z) = (`AO26HSX05_D_F_Z_R,`AO26HSX05_D_R_Z_F);
      (C -=> Z) = (`AO26HSX05_C_F_Z_R,`AO26HSX05_C_R_Z_F);
      (B -=> Z) = (`AO26HSX05_B_F_Z_R,`AO26HSX05_B_R_Z_F);
      (A -=> Z) = (`AO26HSX05_A_F_Z_R,`AO26HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // AO26HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:08:53 and Version :1.1 //
 
//  START 
// CELL AO26NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO26NHS_E_F_Z_F 0.1
`define AO26NHS_E_R_Z_R 0.1
`define AO26NHS_D_F_Z_F 0.1
`define AO26NHS_D_R_Z_R 0.1
`define AO26NHS_C_F_Z_F 0.1
`define AO26NHS_C_R_Z_R 0.1
`define AO26NHS_B_F_Z_F 0.1
`define AO26NHS_B_R_Z_R 0.1
`define AO26NHS_A_F_Z_F 0.1
`define AO26NHS_A_R_Z_R 0.1

module AO26NHS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndAB_, A, B);
   or  u1 (OrAndAB_CD_, AndAB_, C, D);
   and  u2 (Z, OrAndAB_CD_, E);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO26NHS_E_R_Z_R,`AO26NHS_E_F_Z_F);
      (D +=> Z) = (`AO26NHS_D_R_Z_R,`AO26NHS_D_F_Z_F);
      (C +=> Z) = (`AO26NHS_C_R_Z_R,`AO26NHS_C_F_Z_F);
      (B +=> Z) = (`AO26NHS_B_R_Z_R,`AO26NHS_B_F_Z_F);
      (A +=> Z) = (`AO26NHS_A_R_Z_R,`AO26NHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO26NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:08:23 and Version :1.1 //
 
//  START 
// CELL AO26NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO26NHSP_E_F_Z_F 0.1
`define AO26NHSP_E_R_Z_R 0.1
`define AO26NHSP_D_F_Z_F 0.1
`define AO26NHSP_D_R_Z_R 0.1
`define AO26NHSP_C_F_Z_F 0.1
`define AO26NHSP_C_R_Z_R 0.1
`define AO26NHSP_B_F_Z_F 0.1
`define AO26NHSP_B_R_Z_R 0.1
`define AO26NHSP_A_F_Z_F 0.1
`define AO26NHSP_A_R_Z_R 0.1

module AO26NHSP (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndAB_, A, B);
   or  u1 (OrAndAB_CD_, AndAB_, C, D);
   and  u2 (Z, OrAndAB_CD_, E);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO26NHSP_E_R_Z_R,`AO26NHSP_E_F_Z_F);
      (D +=> Z) = (`AO26NHSP_D_R_Z_R,`AO26NHSP_D_F_Z_F);
      (C +=> Z) = (`AO26NHSP_C_R_Z_R,`AO26NHSP_C_F_Z_F);
      (B +=> Z) = (`AO26NHSP_B_R_Z_R,`AO26NHSP_B_F_Z_F);
      (A +=> Z) = (`AO26NHSP_A_R_Z_R,`AO26NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO26NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:08:23 and Version :1.1 //
 
//  START 
// CELL AO27HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO27HSX05_E_F_Z_R 0.1
`define AO27HSX05_E_R_Z_F 0.1
`define AO27HSX05_D_F_Z_R 0.1
`define AO27HSX05_D_R_Z_F 0.1
`define AO27HSX05_C_F_Z_R 0.1
`define AO27HSX05_C_R_Z_F 0.1
`define AO27HSX05_B_F_Z_R 0.1
`define AO27HSX05_B_R_Z_F 0.1
`define AO27HSX05_A_F_Z_R 0.1
`define AO27HSX05_A_R_Z_F 0.1

module AO27HSX05 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndABD_, A, B, D);
   and  u1 (AndCD_, C, D);
   nor  u2 (Z, AndABD_, E, AndCD_);


`ifdef functional
`else
   specify

      (E -=> Z) = (`AO27HSX05_E_F_Z_R,`AO27HSX05_E_R_Z_F);
      (D -=> Z) = (`AO27HSX05_D_F_Z_R,`AO27HSX05_D_R_Z_F);
      (C -=> Z) = (`AO27HSX05_C_F_Z_R,`AO27HSX05_C_R_Z_F);
      (B -=> Z) = (`AO27HSX05_B_F_Z_R,`AO27HSX05_B_R_Z_F);
      (A -=> Z) = (`AO27HSX05_A_F_Z_R,`AO27HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // AO27HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:04 and Version :1.1 //
 
//  START 
// CELL AO27NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO27NHS_E_F_Z_F 0.1
`define AO27NHS_E_R_Z_R 0.1
`define AO27NHS_D_F_Z_F 0.1
`define AO27NHS_D_R_Z_R 0.1
`define AO27NHS_C_F_Z_F 0.1
`define AO27NHS_C_R_Z_R 0.1
`define AO27NHS_B_F_Z_F 0.1
`define AO27NHS_B_R_Z_R 0.1
`define AO27NHS_A_F_Z_F 0.1
`define AO27NHS_A_R_Z_R 0.1

module AO27NHS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndABD_, A, B, D);
   and  u1 (AndCD_, C, D);
   or  u2 (Z, AndABD_, E, AndCD_);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO27NHS_E_R_Z_R,`AO27NHS_E_F_Z_F);
      (D +=> Z) = (`AO27NHS_D_R_Z_R,`AO27NHS_D_F_Z_F);
      (C +=> Z) = (`AO27NHS_C_R_Z_R,`AO27NHS_C_F_Z_F);
      (B +=> Z) = (`AO27NHS_B_R_Z_R,`AO27NHS_B_F_Z_F);
      (A +=> Z) = (`AO27NHS_A_R_Z_R,`AO27NHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO27NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:08:53 and Version :1.1 //
 
//  START 
// CELL AO27NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO27NHSP_E_F_Z_F 0.1
`define AO27NHSP_E_R_Z_R 0.1
`define AO27NHSP_D_F_Z_F 0.1
`define AO27NHSP_D_R_Z_R 0.1
`define AO27NHSP_C_F_Z_F 0.1
`define AO27NHSP_C_R_Z_R 0.1
`define AO27NHSP_B_F_Z_F 0.1
`define AO27NHSP_B_R_Z_R 0.1
`define AO27NHSP_A_F_Z_F 0.1
`define AO27NHSP_A_R_Z_R 0.1

module AO27NHSP (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndABD_, A, B, D);
   and  u1 (AndCD_, C, D);
   or  u2 (Z, AndABD_, E, AndCD_);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO27NHSP_E_R_Z_R,`AO27NHSP_E_F_Z_F);
      (D +=> Z) = (`AO27NHSP_D_R_Z_R,`AO27NHSP_D_F_Z_F);
      (C +=> Z) = (`AO27NHSP_C_R_Z_R,`AO27NHSP_C_F_Z_F);
      (B +=> Z) = (`AO27NHSP_B_R_Z_R,`AO27NHSP_B_F_Z_F);
      (A +=> Z) = (`AO27NHSP_A_R_Z_R,`AO27NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO27NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:08:53 and Version :1.1 //
 
//  START 
// CELL AO2AHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO2AHS_D_F_Z_R 0.1
`define AO2AHS_D_R_Z_F 0.1
`define AO2AHS_C_F_Z_R 0.1
`define AO2AHS_C_R_Z_F 0.1
`define AO2AHS_B_F_Z_R 0.1
`define AO2AHS_B_R_Z_F 0.1
`define AO2AHS_A_F_Z_F 0.1
`define AO2AHS_A_R_Z_R 0.1

module AO2AHS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAXB_, AndCD_);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAXB_, AX, B);
   not  u3 (AX, A);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO2AHS_D_F_Z_R,`AO2AHS_D_R_Z_F);
      (C -=> Z) = (`AO2AHS_C_F_Z_R,`AO2AHS_C_R_Z_F);
      (B -=> Z) = (`AO2AHS_B_F_Z_R,`AO2AHS_B_R_Z_F);
      (A +=> Z) = (`AO2AHS_A_R_Z_R,`AO2AHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO2AHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:07 and Version :1.1 //
 
//  START 
// CELL AO2AHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO2AHSP_D_F_Z_R 0.1
`define AO2AHSP_D_R_Z_F 0.1
`define AO2AHSP_C_F_Z_R 0.1
`define AO2AHSP_C_R_Z_F 0.1
`define AO2AHSP_B_F_Z_R 0.1
`define AO2AHSP_B_R_Z_F 0.1
`define AO2AHSP_A_F_Z_F 0.1
`define AO2AHSP_A_R_Z_R 0.1

module AO2AHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAXB_, AndCD_);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAXB_, AX, B);
   not  u3 (AX, A);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO2AHSP_D_F_Z_R,`AO2AHSP_D_R_Z_F);
      (C -=> Z) = (`AO2AHSP_C_F_Z_R,`AO2AHSP_C_R_Z_F);
      (B -=> Z) = (`AO2AHSP_B_F_Z_R,`AO2AHSP_B_R_Z_F);
      (A +=> Z) = (`AO2AHSP_A_R_Z_R,`AO2AHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO2AHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:07 and Version :1.1 //
 
//  START 
// CELL AO2AHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO2AHSX4_D_F_Z_R 0.1
`define AO2AHSX4_D_R_Z_F 0.1
`define AO2AHSX4_C_F_Z_R 0.1
`define AO2AHSX4_C_R_Z_F 0.1
`define AO2AHSX4_B_F_Z_R 0.1
`define AO2AHSX4_B_R_Z_F 0.1
`define AO2AHSX4_A_F_Z_F 0.1
`define AO2AHSX4_A_R_Z_R 0.1

module AO2AHSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAXB_, AndCD_);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAXB_, AX, B);
   not  u3 (AX, A);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO2AHSX4_D_F_Z_R,`AO2AHSX4_D_R_Z_F);
      (C -=> Z) = (`AO2AHSX4_C_F_Z_R,`AO2AHSX4_C_R_Z_F);
      (B -=> Z) = (`AO2AHSX4_B_F_Z_R,`AO2AHSX4_B_R_Z_F);
      (A +=> Z) = (`AO2AHSX4_A_R_Z_R,`AO2AHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO2AHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:07 and Version :1.1 //
 
//  START 
// CELL AO2AHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO2AHSX8_D_F_Z_R 0.1
`define AO2AHSX8_D_R_Z_F 0.1
`define AO2AHSX8_C_F_Z_R 0.1
`define AO2AHSX8_C_R_Z_F 0.1
`define AO2AHSX8_B_F_Z_R 0.1
`define AO2AHSX8_B_R_Z_F 0.1
`define AO2AHSX8_A_F_Z_F 0.1
`define AO2AHSX8_A_R_Z_R 0.1

module AO2AHSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAXB_, AndCD_);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAXB_, AX, B);
   not  u3 (AX, A);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO2AHSX8_D_F_Z_R,`AO2AHSX8_D_R_Z_F);
      (C -=> Z) = (`AO2AHSX8_C_F_Z_R,`AO2AHSX8_C_R_Z_F);
      (B -=> Z) = (`AO2AHSX8_B_F_Z_R,`AO2AHSX8_B_R_Z_F);
      (A +=> Z) = (`AO2AHSX8_A_R_Z_R,`AO2AHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO2AHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:07 and Version :1.1 //
 
//  START 
// CELL F_AO2AHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO2AHSX4_D_F_Z_R 0.1
`define F_AO2AHSX4_D_R_Z_F 0.1
`define F_AO2AHSX4_C_F_Z_R 0.1
`define F_AO2AHSX4_C_R_Z_F 0.1
`define F_AO2AHSX4_B_F_Z_R 0.1
`define F_AO2AHSX4_B_R_Z_F 0.1
`define F_AO2AHSX4_A_F_Z_F 0.1
`define F_AO2AHSX4_A_R_Z_R 0.1

module F_AO2AHSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, AndAXB_, AndCD_);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAXB_, AX, B);
   not  u3 (AX, A);


`ifdef functional
`else
   specify

      (D -=> Z) = (`F_AO2AHSX4_D_F_Z_R,`F_AO2AHSX4_D_R_Z_F);
      (C -=> Z) = (`F_AO2AHSX4_C_F_Z_R,`F_AO2AHSX4_C_R_Z_F);
      (B -=> Z) = (`F_AO2AHSX4_B_F_Z_R,`F_AO2AHSX4_B_R_Z_F);
      (A +=> Z) = (`F_AO2AHSX4_A_R_Z_R,`F_AO2AHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // F_AO2AHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:07 and Version :1.1 //
 
//  START 
// CELL AO2ANHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO2ANHS_D_F_Z_F 0.1
`define AO2ANHS_D_R_Z_R 0.1
`define AO2ANHS_C_F_Z_F 0.1
`define AO2ANHS_C_R_Z_R 0.1
`define AO2ANHS_B_F_Z_F 0.1
`define AO2ANHS_B_R_Z_R 0.1
`define AO2ANHS_A_F_Z_R 0.1
`define AO2ANHS_A_R_Z_F 0.1

module AO2ANHS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, AndAXB_, AndCD_);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAXB_, AX, B);
   not  u3 (AX, A);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO2ANHS_D_R_Z_R,`AO2ANHS_D_F_Z_F);
      (C +=> Z) = (`AO2ANHS_C_R_Z_R,`AO2ANHS_C_F_Z_F);
      (B +=> Z) = (`AO2ANHS_B_R_Z_R,`AO2ANHS_B_F_Z_F);
      (A -=> Z) = (`AO2ANHS_A_F_Z_R,`AO2ANHS_A_R_Z_F);

   endspecify
`endif


endmodule // AO2ANHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:07 and Version :1.1 //
 
//  START 
// CELL AO2ANHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO2ANHSP_D_F_Z_F 0.1
`define AO2ANHSP_D_R_Z_R 0.1
`define AO2ANHSP_C_F_Z_F 0.1
`define AO2ANHSP_C_R_Z_R 0.1
`define AO2ANHSP_B_F_Z_F 0.1
`define AO2ANHSP_B_R_Z_R 0.1
`define AO2ANHSP_A_F_Z_R 0.1
`define AO2ANHSP_A_R_Z_F 0.1

module AO2ANHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, AndAXB_, AndCD_);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAXB_, AX, B);
   not  u3 (AX, A);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO2ANHSP_D_R_Z_R,`AO2ANHSP_D_F_Z_F);
      (C +=> Z) = (`AO2ANHSP_C_R_Z_R,`AO2ANHSP_C_F_Z_F);
      (B +=> Z) = (`AO2ANHSP_B_R_Z_R,`AO2ANHSP_B_F_Z_F);
      (A -=> Z) = (`AO2ANHSP_A_F_Z_R,`AO2ANHSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO2ANHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:07 and Version :1.1 //
 
//  START 
// CELL AO2ANHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO2ANHSX4_D_F_Z_F 0.1
`define AO2ANHSX4_D_R_Z_R 0.1
`define AO2ANHSX4_C_F_Z_F 0.1
`define AO2ANHSX4_C_R_Z_R 0.1
`define AO2ANHSX4_B_F_Z_F 0.1
`define AO2ANHSX4_B_R_Z_R 0.1
`define AO2ANHSX4_A_F_Z_R 0.1
`define AO2ANHSX4_A_R_Z_F 0.1

module AO2ANHSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, AndAXB_, AndCD_);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAXB_, AX, B);
   not  u3 (AX, A);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO2ANHSX4_D_R_Z_R,`AO2ANHSX4_D_F_Z_F);
      (C +=> Z) = (`AO2ANHSX4_C_R_Z_R,`AO2ANHSX4_C_F_Z_F);
      (B +=> Z) = (`AO2ANHSX4_B_R_Z_R,`AO2ANHSX4_B_F_Z_F);
      (A -=> Z) = (`AO2ANHSX4_A_F_Z_R,`AO2ANHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO2ANHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:07 and Version :1.1 //
 
//  START 
// CELL AO2ANHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO2ANHSX8_D_F_Z_F 0.1
`define AO2ANHSX8_D_R_Z_R 0.1
`define AO2ANHSX8_C_F_Z_F 0.1
`define AO2ANHSX8_C_R_Z_R 0.1
`define AO2ANHSX8_B_F_Z_F 0.1
`define AO2ANHSX8_B_R_Z_R 0.1
`define AO2ANHSX8_A_F_Z_R 0.1
`define AO2ANHSX8_A_R_Z_F 0.1

module AO2ANHSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, AndAXB_, AndCD_);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAXB_, AX, B);
   not  u3 (AX, A);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO2ANHSX8_D_R_Z_R,`AO2ANHSX8_D_F_Z_F);
      (C +=> Z) = (`AO2ANHSX8_C_R_Z_R,`AO2ANHSX8_C_F_Z_F);
      (B +=> Z) = (`AO2ANHSX8_B_R_Z_R,`AO2ANHSX8_B_F_Z_F);
      (A -=> Z) = (`AO2ANHSX8_A_F_Z_R,`AO2ANHSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AO2ANHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:07 and Version :1.1 //
 
//  START 
// CELL AO2NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO2NHS_D_F_Z_F 0.1
`define AO2NHS_D_R_Z_R 0.1
`define AO2NHS_C_F_Z_F 0.1
`define AO2NHS_C_R_Z_R 0.1
`define AO2NHS_B_F_Z_F 0.1
`define AO2NHS_B_R_Z_R 0.1
`define AO2NHS_A_F_Z_F 0.1
`define AO2NHS_A_R_Z_R 0.1

module AO2NHS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, AndAB_, AndCD_);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO2NHS_D_R_Z_R,`AO2NHS_D_F_Z_F);
      (C +=> Z) = (`AO2NHS_C_R_Z_R,`AO2NHS_C_F_Z_F);
      (B +=> Z) = (`AO2NHS_B_R_Z_R,`AO2NHS_B_F_Z_F);
      (A +=> Z) = (`AO2NHS_A_R_Z_R,`AO2NHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO2NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:09 and Version :1.1 //
 
//  START 
// CELL AO2NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO2NHSP_D_F_Z_F 0.1
`define AO2NHSP_D_R_Z_R 0.1
`define AO2NHSP_C_F_Z_F 0.1
`define AO2NHSP_C_R_Z_R 0.1
`define AO2NHSP_B_F_Z_F 0.1
`define AO2NHSP_B_R_Z_R 0.1
`define AO2NHSP_A_F_Z_F 0.1
`define AO2NHSP_A_R_Z_R 0.1

module AO2NHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, AndAB_, AndCD_);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO2NHSP_D_R_Z_R,`AO2NHSP_D_F_Z_F);
      (C +=> Z) = (`AO2NHSP_C_R_Z_R,`AO2NHSP_C_F_Z_F);
      (B +=> Z) = (`AO2NHSP_B_R_Z_R,`AO2NHSP_B_F_Z_F);
      (A +=> Z) = (`AO2NHSP_A_R_Z_R,`AO2NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO2NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:09 and Version :1.1 //
 
//  START 
// CELL AO2NHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO2NHSX4_D_F_Z_F 0.1
`define AO2NHSX4_D_R_Z_R 0.1
`define AO2NHSX4_C_F_Z_F 0.1
`define AO2NHSX4_C_R_Z_R 0.1
`define AO2NHSX4_B_F_Z_F 0.1
`define AO2NHSX4_B_R_Z_R 0.1
`define AO2NHSX4_A_F_Z_F 0.1
`define AO2NHSX4_A_R_Z_R 0.1

module AO2NHSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, AndAB_, AndCD_);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO2NHSX4_D_R_Z_R,`AO2NHSX4_D_F_Z_F);
      (C +=> Z) = (`AO2NHSX4_C_R_Z_R,`AO2NHSX4_C_F_Z_F);
      (B +=> Z) = (`AO2NHSX4_B_R_Z_R,`AO2NHSX4_B_F_Z_F);
      (A +=> Z) = (`AO2NHSX4_A_R_Z_R,`AO2NHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO2NHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:09 and Version :1.1 //
 
//  START 
// CELL AO2NHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO2NHSX8_D_F_Z_F 0.1
`define AO2NHSX8_D_R_Z_R 0.1
`define AO2NHSX8_C_F_Z_F 0.1
`define AO2NHSX8_C_R_Z_R 0.1
`define AO2NHSX8_B_F_Z_F 0.1
`define AO2NHSX8_B_R_Z_R 0.1
`define AO2NHSX8_A_F_Z_F 0.1
`define AO2NHSX8_A_R_Z_R 0.1

module AO2NHSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, AndAB_, AndCD_);
   and  u1 (AndCD_, C, D);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO2NHSX8_D_R_Z_R,`AO2NHSX8_D_F_Z_F);
      (C +=> Z) = (`AO2NHSX8_C_R_Z_R,`AO2NHSX8_C_F_Z_F);
      (B +=> Z) = (`AO2NHSX8_B_R_Z_R,`AO2NHSX8_B_F_Z_F);
      (A +=> Z) = (`AO2NHSX8_A_R_Z_R,`AO2NHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO2NHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:09 and Version :1.1 //
 
//  START 
// CELL AO3HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3HSX05_D_F_Z_R 0.1
`define AO3HSX05_D_R_Z_F 0.1
`define AO3HSX05_C_F_Z_R 0.1
`define AO3HSX05_C_R_Z_F 0.1
`define AO3HSX05_B_F_Z_R 0.1
`define AO3HSX05_B_R_Z_F 0.1
`define AO3HSX05_A_F_Z_R 0.1
`define AO3HSX05_A_R_Z_F 0.1

module AO3HSX05 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAB_, C, D);
   or  u1 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO3HSX05_D_F_Z_R,`AO3HSX05_D_R_Z_F);
      (C -=> Z) = (`AO3HSX05_C_F_Z_R,`AO3HSX05_C_R_Z_F);
      (B -=> Z) = (`AO3HSX05_B_F_Z_R,`AO3HSX05_B_R_Z_F);
      (A -=> Z) = (`AO3HSX05_A_F_Z_R,`AO3HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // AO3HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:45 and Version :1.1 //
 
//  START 
// CELL AO3HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3HS_D_F_Z_R 0.1
`define AO3HS_D_R_Z_F 0.1
`define AO3HS_C_F_Z_R 0.1
`define AO3HS_C_R_Z_F 0.1
`define AO3HS_B_F_Z_R 0.1
`define AO3HS_B_R_Z_F 0.1
`define AO3HS_A_F_Z_R 0.1
`define AO3HS_A_R_Z_F 0.1

module AO3HS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAB_, C, D);
   or  u1 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO3HS_D_F_Z_R,`AO3HS_D_R_Z_F);
      (C -=> Z) = (`AO3HS_C_F_Z_R,`AO3HS_C_R_Z_F);
      (B -=> Z) = (`AO3HS_B_F_Z_R,`AO3HS_B_R_Z_F);
      (A -=> Z) = (`AO3HS_A_F_Z_R,`AO3HS_A_R_Z_F);

   endspecify
`endif


endmodule // AO3HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:45 and Version :1.1 //
 
//  START 
// CELL AO3HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3HSP_D_F_Z_R 0.1
`define AO3HSP_D_R_Z_F 0.1
`define AO3HSP_C_F_Z_R 0.1
`define AO3HSP_C_R_Z_F 0.1
`define AO3HSP_B_F_Z_R 0.1
`define AO3HSP_B_R_Z_F 0.1
`define AO3HSP_A_F_Z_R 0.1
`define AO3HSP_A_R_Z_F 0.1

module AO3HSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAB_, C, D);
   or  u1 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO3HSP_D_F_Z_R,`AO3HSP_D_R_Z_F);
      (C -=> Z) = (`AO3HSP_C_F_Z_R,`AO3HSP_C_R_Z_F);
      (B -=> Z) = (`AO3HSP_B_F_Z_R,`AO3HSP_B_R_Z_F);
      (A -=> Z) = (`AO3HSP_A_F_Z_R,`AO3HSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO3HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:45 and Version :1.1 //
 
//  START 
// CELL AO3HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3HSX4_D_F_Z_R 0.1
`define AO3HSX4_D_R_Z_F 0.1
`define AO3HSX4_C_F_Z_R 0.1
`define AO3HSX4_C_R_Z_F 0.1
`define AO3HSX4_B_F_Z_R 0.1
`define AO3HSX4_B_R_Z_F 0.1
`define AO3HSX4_A_F_Z_R 0.1
`define AO3HSX4_A_R_Z_F 0.1

module AO3HSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAB_, C, D);
   or  u1 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO3HSX4_D_F_Z_R,`AO3HSX4_D_R_Z_F);
      (C -=> Z) = (`AO3HSX4_C_F_Z_R,`AO3HSX4_C_R_Z_F);
      (B -=> Z) = (`AO3HSX4_B_F_Z_R,`AO3HSX4_B_R_Z_F);
      (A -=> Z) = (`AO3HSX4_A_F_Z_R,`AO3HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO3HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:45 and Version :1.1 //
 
//  START 
// CELL AO3HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3HSX8_D_F_Z_R 0.1
`define AO3HSX8_D_R_Z_F 0.1
`define AO3HSX8_C_F_Z_R 0.1
`define AO3HSX8_C_R_Z_F 0.1
`define AO3HSX8_B_F_Z_R 0.1
`define AO3HSX8_B_R_Z_F 0.1
`define AO3HSX8_A_F_Z_R 0.1
`define AO3HSX8_A_R_Z_F 0.1

module AO3HSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAB_, C, D);
   or  u1 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO3HSX8_D_F_Z_R,`AO3HSX8_D_R_Z_F);
      (C -=> Z) = (`AO3HSX8_C_F_Z_R,`AO3HSX8_C_R_Z_F);
      (B -=> Z) = (`AO3HSX8_B_F_Z_R,`AO3HSX8_B_R_Z_F);
      (A -=> Z) = (`AO3HSX8_A_F_Z_R,`AO3HSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AO3HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:45 and Version :1.1 //
 
//  START 
// CELL AO39HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO39HS_F_F_Z_R 0.1
`define AO39HS_F_R_Z_F 0.1
`define AO39HS_E_F_Z_R 0.1
`define AO39HS_E_R_Z_F 0.1
`define AO39HS_D_F_Z_R 0.1
`define AO39HS_D_R_Z_F 0.1
`define AO39HS_C_F_Z_R 0.1
`define AO39HS_C_R_Z_F 0.1
`define AO39HS_B_F_Z_R 0.1
`define AO39HS_B_R_Z_F 0.1
`define AO39HS_A_F_Z_R 0.1
`define AO39HS_A_R_Z_F 0.1

module AO39HS (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   nand  u0 (Z, OrAB_, OrCD_, OrEF_);
   or  u1 (OrEF_, E, F);
   or  u2 (OrCD_, C, D);
   or  u3 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (F -=> Z) = (`AO39HS_F_F_Z_R,`AO39HS_F_R_Z_F);
      (E -=> Z) = (`AO39HS_E_F_Z_R,`AO39HS_E_R_Z_F);
      (D -=> Z) = (`AO39HS_D_F_Z_R,`AO39HS_D_R_Z_F);
      (C -=> Z) = (`AO39HS_C_F_Z_R,`AO39HS_C_R_Z_F);
      (B -=> Z) = (`AO39HS_B_F_Z_R,`AO39HS_B_R_Z_F);
      (A -=> Z) = (`AO39HS_A_F_Z_R,`AO39HS_A_R_Z_F);

   endspecify
`endif


endmodule // AO39HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:48 and Version :1.1 //
 
//  START 
// CELL F_AO39HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO39HS_F_F_Z_R 0.1
`define F_AO39HS_F_R_Z_F 0.1
`define F_AO39HS_E_F_Z_R 0.1
`define F_AO39HS_E_R_Z_F 0.1
`define F_AO39HS_D_F_Z_R 0.1
`define F_AO39HS_D_R_Z_F 0.1
`define F_AO39HS_C_F_Z_R 0.1
`define F_AO39HS_C_R_Z_F 0.1
`define F_AO39HS_B_F_Z_R 0.1
`define F_AO39HS_B_R_Z_F 0.1
`define F_AO39HS_A_F_Z_R 0.1
`define F_AO39HS_A_R_Z_F 0.1

module F_AO39HS (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   nand  u0 (Z, OrAB_, OrCD_, OrEF_);
   or  u1 (OrEF_, E, F);
   or  u2 (OrCD_, C, D);
   or  u3 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (F -=> Z) = (`F_AO39HS_F_F_Z_R,`F_AO39HS_F_R_Z_F);
      (E -=> Z) = (`F_AO39HS_E_F_Z_R,`F_AO39HS_E_R_Z_F);
      (D -=> Z) = (`F_AO39HS_D_F_Z_R,`F_AO39HS_D_R_Z_F);
      (C -=> Z) = (`F_AO39HS_C_F_Z_R,`F_AO39HS_C_R_Z_F);
      (B -=> Z) = (`F_AO39HS_B_F_Z_R,`F_AO39HS_B_R_Z_F);
      (A -=> Z) = (`F_AO39HS_A_F_Z_R,`F_AO39HS_A_R_Z_F);

   endspecify
`endif


endmodule // F_AO39HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:48 and Version :1.1 //
 
//  START 
// Cell F_AO39NHS 

`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define F_AO39NHS_A_R_Z_R 0.1
`define F_AO39NHS_A_F_Z_F 0.1
`define F_AO39NHS_B_R_Z_R 0.1
`define F_AO39NHS_B_F_Z_F 0.1
`define F_AO39NHS_C_R_Z_R 0.1
`define F_AO39NHS_C_F_Z_F 0.1
`define F_AO39NHS_D_R_Z_R 0.1
`define F_AO39NHS_D_F_Z_F 0.1
`define F_AO39NHS_E_R_Z_R 0.1
`define F_AO39NHS_E_F_Z_F 0.1
`define F_AO39NHS_F_R_Z_R 0.1
`define F_AO39NHS_F_F_Z_F 0.1

module F_AO39NHS  (Z, A, B, C, D, E, F);

	output Z;
	input A;
	input B;
	input C;
	input D;
	input E;
	input F;

	or    U1 (INTERNAL1, A, B) ;
	or    U2 (INTERNAL2, C, D) ;
	or    U3 (INTERNAL3, E, F) ;
	and    U4 (Z, INTERNAL1, INTERNAL2, INTERNAL3) ;


`ifdef functional
`else

	specify

		(A +=> Z) = (`F_AO39NHS_A_R_Z_R,`F_AO39NHS_A_F_Z_F);
		(B +=> Z) = (`F_AO39NHS_B_R_Z_R,`F_AO39NHS_B_F_Z_F);
		(C +=> Z) = (`F_AO39NHS_C_R_Z_R,`F_AO39NHS_C_F_Z_F);
		(D +=> Z) = (`F_AO39NHS_D_R_Z_R,`F_AO39NHS_D_F_Z_F);
		(E +=> Z) = (`F_AO39NHS_E_R_Z_R,`F_AO39NHS_E_F_Z_F);
		(F +=> Z) = (`F_AO39NHS_F_R_Z_R,`F_AO39NHS_F_F_Z_F);


	endspecify

`endif

endmodule // F_AO39NHS

`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine

//  END

// CELL AO3AHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3AHS_D_F_Z_R 0.1
`define AO3AHS_D_R_Z_F 0.1
`define AO3AHS_C_F_Z_R 0.1
`define AO3AHS_C_R_Z_F 0.1
`define AO3AHS_B_F_Z_R 0.1
`define AO3AHS_B_R_Z_F 0.1
`define AO3AHS_A_F_Z_F 0.1
`define AO3AHS_A_R_Z_R 0.1

module AO3AHS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAXB_, C, D);
   or  u1 (OrAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO3AHS_D_F_Z_R,`AO3AHS_D_R_Z_F);
      (C -=> Z) = (`AO3AHS_C_F_Z_R,`AO3AHS_C_R_Z_F);
      (B -=> Z) = (`AO3AHS_B_F_Z_R,`AO3AHS_B_R_Z_F);
      (A +=> Z) = (`AO3AHS_A_R_Z_R,`AO3AHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO3AHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:51 and Version :1.1 //
 
//  START 
// CELL AO3AHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3AHSP_D_F_Z_R 0.1
`define AO3AHSP_D_R_Z_F 0.1
`define AO3AHSP_C_F_Z_R 0.1
`define AO3AHSP_C_R_Z_F 0.1
`define AO3AHSP_B_F_Z_R 0.1
`define AO3AHSP_B_R_Z_F 0.1
`define AO3AHSP_A_F_Z_F 0.1
`define AO3AHSP_A_R_Z_R 0.1

module AO3AHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAXB_, C, D);
   or  u1 (OrAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO3AHSP_D_F_Z_R,`AO3AHSP_D_R_Z_F);
      (C -=> Z) = (`AO3AHSP_C_F_Z_R,`AO3AHSP_C_R_Z_F);
      (B -=> Z) = (`AO3AHSP_B_F_Z_R,`AO3AHSP_B_R_Z_F);
      (A +=> Z) = (`AO3AHSP_A_R_Z_R,`AO3AHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO3AHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:51 and Version :1.1 //
 
//  START 
// CELL AO3AHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3AHSX4_D_F_Z_R 0.1
`define AO3AHSX4_D_R_Z_F 0.1
`define AO3AHSX4_C_F_Z_R 0.1
`define AO3AHSX4_C_R_Z_F 0.1
`define AO3AHSX4_B_F_Z_R 0.1
`define AO3AHSX4_B_R_Z_F 0.1
`define AO3AHSX4_A_F_Z_F 0.1
`define AO3AHSX4_A_R_Z_R 0.1

module AO3AHSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAXB_, C, D);
   or  u1 (OrAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO3AHSX4_D_F_Z_R,`AO3AHSX4_D_R_Z_F);
      (C -=> Z) = (`AO3AHSX4_C_F_Z_R,`AO3AHSX4_C_R_Z_F);
      (B -=> Z) = (`AO3AHSX4_B_F_Z_R,`AO3AHSX4_B_R_Z_F);
      (A +=> Z) = (`AO3AHSX4_A_R_Z_R,`AO3AHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO3AHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:51 and Version :1.1 //
 
//  START 
// CELL AO3AHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3AHSX8_D_F_Z_R 0.1
`define AO3AHSX8_D_R_Z_F 0.1
`define AO3AHSX8_C_F_Z_R 0.1
`define AO3AHSX8_C_R_Z_F 0.1
`define AO3AHSX8_B_F_Z_R 0.1
`define AO3AHSX8_B_R_Z_F 0.1
`define AO3AHSX8_A_F_Z_F 0.1
`define AO3AHSX8_A_R_Z_R 0.1

module AO3AHSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAXB_, C, D);
   or  u1 (OrAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO3AHSX8_D_F_Z_R,`AO3AHSX8_D_R_Z_F);
      (C -=> Z) = (`AO3AHSX8_C_F_Z_R,`AO3AHSX8_C_R_Z_F);
      (B -=> Z) = (`AO3AHSX8_B_F_Z_R,`AO3AHSX8_B_R_Z_F);
      (A +=> Z) = (`AO3AHSX8_A_R_Z_R,`AO3AHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO3AHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:51 and Version :1.1 //
 
//  START 
// CELL F_AO3AHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO3AHSP_D_F_Z_R 0.1
`define F_AO3AHSP_D_R_Z_F 0.1
`define F_AO3AHSP_C_F_Z_R 0.1
`define F_AO3AHSP_C_R_Z_F 0.1
`define F_AO3AHSP_B_F_Z_R 0.1
`define F_AO3AHSP_B_R_Z_F 0.1
`define F_AO3AHSP_A_F_Z_F 0.1
`define F_AO3AHSP_A_R_Z_R 0.1

module F_AO3AHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAXB_, C, D);
   or  u1 (OrAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (D -=> Z) = (`F_AO3AHSP_D_F_Z_R,`F_AO3AHSP_D_R_Z_F);
      (C -=> Z) = (`F_AO3AHSP_C_F_Z_R,`F_AO3AHSP_C_R_Z_F);
      (B -=> Z) = (`F_AO3AHSP_B_F_Z_R,`F_AO3AHSP_B_R_Z_F);
      (A +=> Z) = (`F_AO3AHSP_A_R_Z_R,`F_AO3AHSP_A_F_Z_F);

   endspecify
`endif


endmodule // F_AO3AHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:51 and Version :1.1 //
 
//  START 
// CELL AO3ANHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3ANHS_D_F_Z_F 0.1
`define AO3ANHS_D_R_Z_R 0.1
`define AO3ANHS_C_F_Z_F 0.1
`define AO3ANHS_C_R_Z_R 0.1
`define AO3ANHS_B_F_Z_F 0.1
`define AO3ANHS_B_R_Z_R 0.1
`define AO3ANHS_A_F_Z_R 0.1
`define AO3ANHS_A_R_Z_F 0.1

module AO3ANHS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAXB_, C, D);
   or  u1 (OrAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO3ANHS_D_R_Z_R,`AO3ANHS_D_F_Z_F);
      (C +=> Z) = (`AO3ANHS_C_R_Z_R,`AO3ANHS_C_F_Z_F);
      (B +=> Z) = (`AO3ANHS_B_R_Z_R,`AO3ANHS_B_F_Z_F);
      (A -=> Z) = (`AO3ANHS_A_F_Z_R,`AO3ANHS_A_R_Z_F);

   endspecify
`endif


endmodule // AO3ANHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:51 and Version :1.1 //
 
//  START 
// CELL AO3ANHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3ANHSP_D_F_Z_F 0.1
`define AO3ANHSP_D_R_Z_R 0.1
`define AO3ANHSP_C_F_Z_F 0.1
`define AO3ANHSP_C_R_Z_R 0.1
`define AO3ANHSP_B_F_Z_F 0.1
`define AO3ANHSP_B_R_Z_R 0.1
`define AO3ANHSP_A_F_Z_R 0.1
`define AO3ANHSP_A_R_Z_F 0.1

module AO3ANHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAXB_, C, D);
   or  u1 (OrAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO3ANHSP_D_R_Z_R,`AO3ANHSP_D_F_Z_F);
      (C +=> Z) = (`AO3ANHSP_C_R_Z_R,`AO3ANHSP_C_F_Z_F);
      (B +=> Z) = (`AO3ANHSP_B_R_Z_R,`AO3ANHSP_B_F_Z_F);
      (A -=> Z) = (`AO3ANHSP_A_F_Z_R,`AO3ANHSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO3ANHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:51 and Version :1.1 //
 
//  START 
// CELL AO3ANHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3ANHSX4_D_F_Z_F 0.1
`define AO3ANHSX4_D_R_Z_R 0.1
`define AO3ANHSX4_C_F_Z_F 0.1
`define AO3ANHSX4_C_R_Z_R 0.1
`define AO3ANHSX4_B_F_Z_F 0.1
`define AO3ANHSX4_B_R_Z_R 0.1
`define AO3ANHSX4_A_F_Z_R 0.1
`define AO3ANHSX4_A_R_Z_F 0.1

module AO3ANHSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAXB_, C, D);
   or  u1 (OrAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO3ANHSX4_D_R_Z_R,`AO3ANHSX4_D_F_Z_F);
      (C +=> Z) = (`AO3ANHSX4_C_R_Z_R,`AO3ANHSX4_C_F_Z_F);
      (B +=> Z) = (`AO3ANHSX4_B_R_Z_R,`AO3ANHSX4_B_F_Z_F);
      (A -=> Z) = (`AO3ANHSX4_A_F_Z_R,`AO3ANHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO3ANHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:51 and Version :1.1 //
 
//  START 
// CELL AO3ANHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3ANHSX8_D_F_Z_F 0.1
`define AO3ANHSX8_D_R_Z_R 0.1
`define AO3ANHSX8_C_F_Z_F 0.1
`define AO3ANHSX8_C_R_Z_R 0.1
`define AO3ANHSX8_B_F_Z_F 0.1
`define AO3ANHSX8_B_R_Z_R 0.1
`define AO3ANHSX8_A_F_Z_R 0.1
`define AO3ANHSX8_A_R_Z_F 0.1

module AO3ANHSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAXB_, C, D);
   or  u1 (OrAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO3ANHSX8_D_R_Z_R,`AO3ANHSX8_D_F_Z_F);
      (C +=> Z) = (`AO3ANHSX8_C_R_Z_R,`AO3ANHSX8_C_F_Z_F);
      (B +=> Z) = (`AO3ANHSX8_B_R_Z_R,`AO3ANHSX8_B_F_Z_F);
      (A -=> Z) = (`AO3ANHSX8_A_F_Z_R,`AO3ANHSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AO3ANHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:51 and Version :1.1 //
 
//  START 
// CELL F_AO3ANHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO3ANHSX4_D_F_Z_F 0.1
`define F_AO3ANHSX4_D_R_Z_R 0.1
`define F_AO3ANHSX4_C_F_Z_F 0.1
`define F_AO3ANHSX4_C_R_Z_R 0.1
`define F_AO3ANHSX4_B_F_Z_F 0.1
`define F_AO3ANHSX4_B_R_Z_R 0.1
`define F_AO3ANHSX4_A_F_Z_R 0.1
`define F_AO3ANHSX4_A_R_Z_F 0.1

module F_AO3ANHSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAXB_, C, D);
   or  u1 (OrAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (D +=> Z) = (`F_AO3ANHSX4_D_R_Z_R,`F_AO3ANHSX4_D_F_Z_F);
      (C +=> Z) = (`F_AO3ANHSX4_C_R_Z_R,`F_AO3ANHSX4_C_F_Z_F);
      (B +=> Z) = (`F_AO3ANHSX4_B_R_Z_R,`F_AO3ANHSX4_B_F_Z_F);
      (A -=> Z) = (`F_AO3ANHSX4_A_F_Z_R,`F_AO3ANHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // F_AO3ANHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:51 and Version :1.1 //
 
//  START 
// CELL AO3CHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3CHS_D_F_Z_R 0.1
`define AO3CHS_D_R_Z_F 0.1
`define AO3CHS_C_F_Z_F 0.1
`define AO3CHS_C_R_Z_R 0.1
`define AO3CHS_B_F_Z_R 0.1
`define AO3CHS_B_R_Z_F 0.1
`define AO3CHS_A_F_Z_R 0.1
`define AO3CHS_A_R_Z_F 0.1

module AO3CHS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAB_, CX, D);
   not  u1 (CX, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO3CHS_D_F_Z_R,`AO3CHS_D_R_Z_F);
      (C +=> Z) = (`AO3CHS_C_R_Z_R,`AO3CHS_C_F_Z_F);
      (B -=> Z) = (`AO3CHS_B_F_Z_R,`AO3CHS_B_R_Z_F);
      (A -=> Z) = (`AO3CHS_A_F_Z_R,`AO3CHS_A_R_Z_F);

   endspecify
`endif


endmodule // AO3CHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:58 and Version :1.1 //
 
//  START 
// CELL AO3CHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3CHSP_D_F_Z_R 0.1
`define AO3CHSP_D_R_Z_F 0.1
`define AO3CHSP_C_F_Z_F 0.1
`define AO3CHSP_C_R_Z_R 0.1
`define AO3CHSP_B_F_Z_R 0.1
`define AO3CHSP_B_R_Z_F 0.1
`define AO3CHSP_A_F_Z_R 0.1
`define AO3CHSP_A_R_Z_F 0.1

module AO3CHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAB_, CX, D);
   not  u1 (CX, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO3CHSP_D_F_Z_R,`AO3CHSP_D_R_Z_F);
      (C +=> Z) = (`AO3CHSP_C_R_Z_R,`AO3CHSP_C_F_Z_F);
      (B -=> Z) = (`AO3CHSP_B_F_Z_R,`AO3CHSP_B_R_Z_F);
      (A -=> Z) = (`AO3CHSP_A_F_Z_R,`AO3CHSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO3CHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:58 and Version :1.1 //
 
//  START 
// CELL AO3CHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3CHSX4_D_F_Z_R 0.1
`define AO3CHSX4_D_R_Z_F 0.1
`define AO3CHSX4_C_F_Z_F 0.1
`define AO3CHSX4_C_R_Z_R 0.1
`define AO3CHSX4_B_F_Z_R 0.1
`define AO3CHSX4_B_R_Z_F 0.1
`define AO3CHSX4_A_F_Z_R 0.1
`define AO3CHSX4_A_R_Z_F 0.1

module AO3CHSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAB_, CX, D);
   not  u1 (CX, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO3CHSX4_D_F_Z_R,`AO3CHSX4_D_R_Z_F);
      (C +=> Z) = (`AO3CHSX4_C_R_Z_R,`AO3CHSX4_C_F_Z_F);
      (B -=> Z) = (`AO3CHSX4_B_F_Z_R,`AO3CHSX4_B_R_Z_F);
      (A -=> Z) = (`AO3CHSX4_A_F_Z_R,`AO3CHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO3CHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:58 and Version :1.1 //
 
//  START 
// CELL AO3CHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3CHSX8_D_F_Z_R 0.1
`define AO3CHSX8_D_R_Z_F 0.1
`define AO3CHSX8_C_F_Z_F 0.1
`define AO3CHSX8_C_R_Z_R 0.1
`define AO3CHSX8_B_F_Z_R 0.1
`define AO3CHSX8_B_R_Z_F 0.1
`define AO3CHSX8_A_F_Z_R 0.1
`define AO3CHSX8_A_R_Z_F 0.1

module AO3CHSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAB_, CX, D);
   not  u1 (CX, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO3CHSX8_D_F_Z_R,`AO3CHSX8_D_R_Z_F);
      (C +=> Z) = (`AO3CHSX8_C_R_Z_R,`AO3CHSX8_C_F_Z_F);
      (B -=> Z) = (`AO3CHSX8_B_F_Z_R,`AO3CHSX8_B_R_Z_F);
      (A -=> Z) = (`AO3CHSX8_A_F_Z_R,`AO3CHSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AO3CHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:58 and Version :1.1 //
 
//  START 
// CELL F_AO3CHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO3CHSP_D_F_Z_R 0.1
`define F_AO3CHSP_D_R_Z_F 0.1
`define F_AO3CHSP_C_F_Z_F 0.1
`define F_AO3CHSP_C_R_Z_R 0.1
`define F_AO3CHSP_B_F_Z_R 0.1
`define F_AO3CHSP_B_R_Z_F 0.1
`define F_AO3CHSP_A_F_Z_R 0.1
`define F_AO3CHSP_A_R_Z_F 0.1

module F_AO3CHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAB_, CX, D);
   not  u1 (CX, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`F_AO3CHSP_D_F_Z_R,`F_AO3CHSP_D_R_Z_F);
      (C +=> Z) = (`F_AO3CHSP_C_R_Z_R,`F_AO3CHSP_C_F_Z_F);
      (B -=> Z) = (`F_AO3CHSP_B_F_Z_R,`F_AO3CHSP_B_R_Z_F);
      (A -=> Z) = (`F_AO3CHSP_A_F_Z_R,`F_AO3CHSP_A_R_Z_F);

   endspecify
`endif


endmodule // F_AO3CHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:58 and Version :1.1 //
 
//  START 
// CELL AO3CNHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3CNHS_D_F_Z_F 0.1
`define AO3CNHS_D_R_Z_R 0.1
`define AO3CNHS_C_F_Z_R 0.1
`define AO3CNHS_C_R_Z_F 0.1
`define AO3CNHS_B_F_Z_F 0.1
`define AO3CNHS_B_R_Z_R 0.1
`define AO3CNHS_A_F_Z_F 0.1
`define AO3CNHS_A_R_Z_R 0.1

module AO3CNHS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAB_, CX, D);
   not  u1 (CX, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO3CNHS_D_R_Z_R,`AO3CNHS_D_F_Z_F);
      (C -=> Z) = (`AO3CNHS_C_F_Z_R,`AO3CNHS_C_R_Z_F);
      (B +=> Z) = (`AO3CNHS_B_R_Z_R,`AO3CNHS_B_F_Z_F);
      (A +=> Z) = (`AO3CNHS_A_R_Z_R,`AO3CNHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO3CNHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:58 and Version :1.1 //
 
//  START 
// CELL AO3CNHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3CNHSP_D_F_Z_F 0.1
`define AO3CNHSP_D_R_Z_R 0.1
`define AO3CNHSP_C_F_Z_R 0.1
`define AO3CNHSP_C_R_Z_F 0.1
`define AO3CNHSP_B_F_Z_F 0.1
`define AO3CNHSP_B_R_Z_R 0.1
`define AO3CNHSP_A_F_Z_F 0.1
`define AO3CNHSP_A_R_Z_R 0.1

module AO3CNHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAB_, CX, D);
   not  u1 (CX, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO3CNHSP_D_R_Z_R,`AO3CNHSP_D_F_Z_F);
      (C -=> Z) = (`AO3CNHSP_C_F_Z_R,`AO3CNHSP_C_R_Z_F);
      (B +=> Z) = (`AO3CNHSP_B_R_Z_R,`AO3CNHSP_B_F_Z_F);
      (A +=> Z) = (`AO3CNHSP_A_R_Z_R,`AO3CNHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO3CNHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:58 and Version :1.1 //
 
//  START 
// CELL AO3CNHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3CNHSX4_D_F_Z_F 0.1
`define AO3CNHSX4_D_R_Z_R 0.1
`define AO3CNHSX4_C_F_Z_R 0.1
`define AO3CNHSX4_C_R_Z_F 0.1
`define AO3CNHSX4_B_F_Z_F 0.1
`define AO3CNHSX4_B_R_Z_R 0.1
`define AO3CNHSX4_A_F_Z_F 0.1
`define AO3CNHSX4_A_R_Z_R 0.1

module AO3CNHSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAB_, CX, D);
   not  u1 (CX, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO3CNHSX4_D_R_Z_R,`AO3CNHSX4_D_F_Z_F);
      (C -=> Z) = (`AO3CNHSX4_C_F_Z_R,`AO3CNHSX4_C_R_Z_F);
      (B +=> Z) = (`AO3CNHSX4_B_R_Z_R,`AO3CNHSX4_B_F_Z_F);
      (A +=> Z) = (`AO3CNHSX4_A_R_Z_R,`AO3CNHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO3CNHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:58 and Version :1.1 //
 
//  START 
// CELL AO3CNHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3CNHSX8_D_F_Z_F 0.1
`define AO3CNHSX8_D_R_Z_R 0.1
`define AO3CNHSX8_C_F_Z_R 0.1
`define AO3CNHSX8_C_R_Z_F 0.1
`define AO3CNHSX8_B_F_Z_F 0.1
`define AO3CNHSX8_B_R_Z_R 0.1
`define AO3CNHSX8_A_F_Z_F 0.1
`define AO3CNHSX8_A_R_Z_R 0.1

module AO3CNHSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAB_, CX, D);
   not  u1 (CX, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO3CNHSX8_D_R_Z_R,`AO3CNHSX8_D_F_Z_F);
      (C -=> Z) = (`AO3CNHSX8_C_F_Z_R,`AO3CNHSX8_C_R_Z_F);
      (B +=> Z) = (`AO3CNHSX8_B_R_Z_R,`AO3CNHSX8_B_F_Z_F);
      (A +=> Z) = (`AO3CNHSX8_A_R_Z_R,`AO3CNHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO3CNHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:09:58 and Version :1.1 //
 
//  START 
// CELL AO3NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3NHS_D_F_Z_F 0.1
`define AO3NHS_D_R_Z_R 0.1
`define AO3NHS_C_F_Z_F 0.1
`define AO3NHS_C_R_Z_R 0.1
`define AO3NHS_B_F_Z_F 0.1
`define AO3NHS_B_R_Z_R 0.1
`define AO3NHS_A_F_Z_F 0.1
`define AO3NHS_A_R_Z_R 0.1

module AO3NHS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAB_, C, D);
   or  u1 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO3NHS_D_R_Z_R,`AO3NHS_D_F_Z_F);
      (C +=> Z) = (`AO3NHS_C_R_Z_R,`AO3NHS_C_F_Z_F);
      (B +=> Z) = (`AO3NHS_B_R_Z_R,`AO3NHS_B_F_Z_F);
      (A +=> Z) = (`AO3NHS_A_R_Z_R,`AO3NHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO3NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:10:01 and Version :1.1 //
 
//  START 
// CELL AO3NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3NHSP_D_F_Z_F 0.1
`define AO3NHSP_D_R_Z_R 0.1
`define AO3NHSP_C_F_Z_F 0.1
`define AO3NHSP_C_R_Z_R 0.1
`define AO3NHSP_B_F_Z_F 0.1
`define AO3NHSP_B_R_Z_R 0.1
`define AO3NHSP_A_F_Z_F 0.1
`define AO3NHSP_A_R_Z_R 0.1

module AO3NHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAB_, C, D);
   or  u1 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO3NHSP_D_R_Z_R,`AO3NHSP_D_F_Z_F);
      (C +=> Z) = (`AO3NHSP_C_R_Z_R,`AO3NHSP_C_F_Z_F);
      (B +=> Z) = (`AO3NHSP_B_R_Z_R,`AO3NHSP_B_F_Z_F);
      (A +=> Z) = (`AO3NHSP_A_R_Z_R,`AO3NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO3NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:10:01 and Version :1.1 //
 
//  START 
// CELL AO3NHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3NHSX4_D_F_Z_F 0.1
`define AO3NHSX4_D_R_Z_R 0.1
`define AO3NHSX4_C_F_Z_F 0.1
`define AO3NHSX4_C_R_Z_R 0.1
`define AO3NHSX4_B_F_Z_F 0.1
`define AO3NHSX4_B_R_Z_R 0.1
`define AO3NHSX4_A_F_Z_F 0.1
`define AO3NHSX4_A_R_Z_R 0.1

module AO3NHSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAB_, C, D);
   or  u1 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO3NHSX4_D_R_Z_R,`AO3NHSX4_D_F_Z_F);
      (C +=> Z) = (`AO3NHSX4_C_R_Z_R,`AO3NHSX4_C_F_Z_F);
      (B +=> Z) = (`AO3NHSX4_B_R_Z_R,`AO3NHSX4_B_F_Z_F);
      (A +=> Z) = (`AO3NHSX4_A_R_Z_R,`AO3NHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO3NHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:10:01 and Version :1.1 //
 
//  START 
// CELL AO3NHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO3NHSX8_D_F_Z_F 0.1
`define AO3NHSX8_D_R_Z_R 0.1
`define AO3NHSX8_C_F_Z_F 0.1
`define AO3NHSX8_C_R_Z_R 0.1
`define AO3NHSX8_B_F_Z_F 0.1
`define AO3NHSX8_B_R_Z_R 0.1
`define AO3NHSX8_A_F_Z_F 0.1
`define AO3NHSX8_A_R_Z_R 0.1

module AO3NHSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAB_, C, D);
   or  u1 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO3NHSX8_D_R_Z_R,`AO3NHSX8_D_F_Z_F);
      (C +=> Z) = (`AO3NHSX8_C_R_Z_R,`AO3NHSX8_C_F_Z_F);
      (B +=> Z) = (`AO3NHSX8_B_R_Z_R,`AO3NHSX8_B_F_Z_F);
      (A +=> Z) = (`AO3NHSX8_A_R_Z_R,`AO3NHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO3NHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:10:01 and Version :1.1 //
 
//  START 
// CELL AO4HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO4HSX05_D_F_Z_R 0.1
`define AO4HSX05_D_R_Z_F 0.1
`define AO4HSX05_C_F_Z_R 0.1
`define AO4HSX05_C_R_Z_F 0.1
`define AO4HSX05_B_F_Z_R 0.1
`define AO4HSX05_B_R_Z_F 0.1
`define AO4HSX05_A_F_Z_R 0.1
`define AO4HSX05_A_R_Z_F 0.1

module AO4HSX05 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAB_, OrCD_);
   or  u1 (OrCD_, C, D);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO4HSX05_D_F_Z_R,`AO4HSX05_D_R_Z_F);
      (C -=> Z) = (`AO4HSX05_C_F_Z_R,`AO4HSX05_C_R_Z_F);
      (B -=> Z) = (`AO4HSX05_B_F_Z_R,`AO4HSX05_B_R_Z_F);
      (A -=> Z) = (`AO4HSX05_A_F_Z_R,`AO4HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // AO4HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:10:07 and Version :1.1 //
 
//  START 
// CELL AO4HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO4HS_D_F_Z_R 0.1
`define AO4HS_D_R_Z_F 0.1
`define AO4HS_C_F_Z_R 0.1
`define AO4HS_C_R_Z_F 0.1
`define AO4HS_B_F_Z_R 0.1
`define AO4HS_B_R_Z_F 0.1
`define AO4HS_A_F_Z_R 0.1
`define AO4HS_A_R_Z_F 0.1

module AO4HS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAB_, OrCD_);
   or  u1 (OrCD_, C, D);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO4HS_D_F_Z_R,`AO4HS_D_R_Z_F);
      (C -=> Z) = (`AO4HS_C_F_Z_R,`AO4HS_C_R_Z_F);
      (B -=> Z) = (`AO4HS_B_F_Z_R,`AO4HS_B_R_Z_F);
      (A -=> Z) = (`AO4HS_A_F_Z_R,`AO4HS_A_R_Z_F);

   endspecify
`endif


endmodule // AO4HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:10:07 and Version :1.1 //
 
//  START 
// CELL AO4HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO4HSP_D_F_Z_R 0.1
`define AO4HSP_D_R_Z_F 0.1
`define AO4HSP_C_F_Z_R 0.1
`define AO4HSP_C_R_Z_F 0.1
`define AO4HSP_B_F_Z_R 0.1
`define AO4HSP_B_R_Z_F 0.1
`define AO4HSP_A_F_Z_R 0.1
`define AO4HSP_A_R_Z_F 0.1

module AO4HSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAB_, OrCD_);
   or  u1 (OrCD_, C, D);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO4HSP_D_F_Z_R,`AO4HSP_D_R_Z_F);
      (C -=> Z) = (`AO4HSP_C_F_Z_R,`AO4HSP_C_R_Z_F);
      (B -=> Z) = (`AO4HSP_B_F_Z_R,`AO4HSP_B_R_Z_F);
      (A -=> Z) = (`AO4HSP_A_F_Z_R,`AO4HSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO4HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:10:07 and Version :1.1 //
 
//  START 
// CELL AO4HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO4HSX4_D_F_Z_R 0.1
`define AO4HSX4_D_R_Z_F 0.1
`define AO4HSX4_C_F_Z_R 0.1
`define AO4HSX4_C_R_Z_F 0.1
`define AO4HSX4_B_F_Z_R 0.1
`define AO4HSX4_B_R_Z_F 0.1
`define AO4HSX4_A_F_Z_R 0.1
`define AO4HSX4_A_R_Z_F 0.1

module AO4HSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAB_, OrCD_);
   or  u1 (OrCD_, C, D);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO4HSX4_D_F_Z_R,`AO4HSX4_D_R_Z_F);
      (C -=> Z) = (`AO4HSX4_C_F_Z_R,`AO4HSX4_C_R_Z_F);
      (B -=> Z) = (`AO4HSX4_B_F_Z_R,`AO4HSX4_B_R_Z_F);
      (A -=> Z) = (`AO4HSX4_A_F_Z_R,`AO4HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO4HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:10:07 and Version :1.1 //
 
//  START 
// CELL AO4HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO4HSX8_D_F_Z_R 0.1
`define AO4HSX8_D_R_Z_F 0.1
`define AO4HSX8_C_F_Z_R 0.1
`define AO4HSX8_C_R_Z_F 0.1
`define AO4HSX8_B_F_Z_R 0.1
`define AO4HSX8_B_R_Z_F 0.1
`define AO4HSX8_A_F_Z_R 0.1
`define AO4HSX8_A_R_Z_F 0.1

module AO4HSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAB_, OrCD_);
   or  u1 (OrCD_, C, D);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO4HSX8_D_F_Z_R,`AO4HSX8_D_R_Z_F);
      (C -=> Z) = (`AO4HSX8_C_F_Z_R,`AO4HSX8_C_R_Z_F);
      (B -=> Z) = (`AO4HSX8_B_F_Z_R,`AO4HSX8_B_R_Z_F);
      (A -=> Z) = (`AO4HSX8_A_F_Z_R,`AO4HSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AO4HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:10:07 and Version :1.1 //
 
//  START 
// CELL F_AO4HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO4HS_D_F_Z_R 0.1
`define F_AO4HS_D_R_Z_F 0.1
`define F_AO4HS_C_F_Z_R 0.1
`define F_AO4HS_C_R_Z_F 0.1
`define F_AO4HS_B_F_Z_R 0.1
`define F_AO4HS_B_R_Z_F 0.1
`define F_AO4HS_A_F_Z_R 0.1
`define F_AO4HS_A_R_Z_F 0.1

module F_AO4HS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAB_, OrCD_);
   or  u1 (OrCD_, C, D);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D -=> Z) = (`F_AO4HS_D_F_Z_R,`F_AO4HS_D_R_Z_F);
      (C -=> Z) = (`F_AO4HS_C_F_Z_R,`F_AO4HS_C_R_Z_F);
      (B -=> Z) = (`F_AO4HS_B_F_Z_R,`F_AO4HS_B_R_Z_F);
      (A -=> Z) = (`F_AO4HS_A_F_Z_R,`F_AO4HS_A_R_Z_F);

   endspecify
`endif


endmodule // F_AO4HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:10:07 and Version :1.1 //
 
//  START 
// CELL AO40HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO40HS_D_F_Z_F 0.1
`define AO40HS_D_R_Z_R 0.1
`define AO40HS_C_F_Z_F 0.1
`define AO40HS_C_R_Z_R 0.1
`define AO40HS_B_F_Z_R 0.1
`define AO40HS_B_R_Z_F 0.1
`define AO40HS_A_F_Z_R 0.1
`define AO40HS_A_R_Z_F 0.1

module AO40HS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAXBX_, OrCD_);
   or  u1 (OrCD_, C, D);
   or  u2 (OrAXBX_, AX, BX);
   not  u3 (BX, B);
   not  u4 (AX, A);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO40HS_D_R_Z_R,`AO40HS_D_F_Z_F);
      (C +=> Z) = (`AO40HS_C_R_Z_R,`AO40HS_C_F_Z_F);
      (B -=> Z) = (`AO40HS_B_F_Z_R,`AO40HS_B_R_Z_F);
      (A -=> Z) = (`AO40HS_A_F_Z_R,`AO40HS_A_R_Z_F);

   endspecify
`endif


endmodule // AO40HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:10:07 and Version :1.1 //
 
//  START 
// CELL AO40HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO40HSP_D_F_Z_F 0.1
`define AO40HSP_D_R_Z_R 0.1
`define AO40HSP_C_F_Z_F 0.1
`define AO40HSP_C_R_Z_R 0.1
`define AO40HSP_B_F_Z_R 0.1
`define AO40HSP_B_R_Z_F 0.1
`define AO40HSP_A_F_Z_R 0.1
`define AO40HSP_A_R_Z_F 0.1

module AO40HSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAXBX_, OrCD_);
   or  u1 (OrCD_, C, D);
   or  u2 (OrAXBX_, AX, BX);
   not  u3 (BX, B);
   not  u4 (AX, A);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO40HSP_D_R_Z_R,`AO40HSP_D_F_Z_F);
      (C +=> Z) = (`AO40HSP_C_R_Z_R,`AO40HSP_C_F_Z_F);
      (B -=> Z) = (`AO40HSP_B_F_Z_R,`AO40HSP_B_R_Z_F);
      (A -=> Z) = (`AO40HSP_A_F_Z_R,`AO40HSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO40HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:10:07 and Version :1.1 //
 
//  START 
// CELL AO41HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO41HS_D_F_Z_F 0.1
`define AO41HS_D_R_Z_R 0.1
`define AO41HS_C_F_Z_F 0.1
`define AO41HS_C_R_Z_R 0.1
`define AO41HS_B_F_Z_R 0.1
`define AO41HS_B_R_Z_F 0.1
`define AO41HS_A_F_Z_R 0.1
`define AO41HS_A_R_Z_F 0.1

module AO41HS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, AX, BX, C, D);
   not  u1 (BX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO41HS_D_R_Z_R,`AO41HS_D_F_Z_F);
      (C +=> Z) = (`AO41HS_C_R_Z_R,`AO41HS_C_F_Z_F);
      (B -=> Z) = (`AO41HS_B_F_Z_R,`AO41HS_B_R_Z_F);
      (A -=> Z) = (`AO41HS_A_F_Z_R,`AO41HS_A_R_Z_F);

   endspecify
`endif


endmodule // AO41HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:10:09 and Version :1.1 //
 
//  START 
// CELL AO41HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO41HSP_D_F_Z_F 0.1
`define AO41HSP_D_R_Z_R 0.1
`define AO41HSP_C_F_Z_F 0.1
`define AO41HSP_C_R_Z_R 0.1
`define AO41HSP_B_F_Z_R 0.1
`define AO41HSP_B_R_Z_F 0.1
`define AO41HSP_A_F_Z_R 0.1
`define AO41HSP_A_R_Z_F 0.1

module AO41HSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, AX, BX, C, D);
   not  u1 (BX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO41HSP_D_R_Z_R,`AO41HSP_D_F_Z_F);
      (C +=> Z) = (`AO41HSP_C_R_Z_R,`AO41HSP_C_F_Z_F);
      (B -=> Z) = (`AO41HSP_B_F_Z_R,`AO41HSP_B_R_Z_F);
      (A -=> Z) = (`AO41HSP_A_F_Z_R,`AO41HSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO41HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:10:09 and Version :1.1 //
 
//  START 
// CELL AO4AHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO4AHS_D_F_Z_R 0.1
`define AO4AHS_D_R_Z_F 0.1
`define AO4AHS_C_F_Z_R 0.1
`define AO4AHS_C_R_Z_F 0.1
`define AO4AHS_B_F_Z_R 0.1
`define AO4AHS_B_R_Z_F 0.1
`define AO4AHS_A_F_Z_F 0.1
`define AO4AHS_A_R_Z_R 0.1

module AO4AHS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAXB_, OrCD_);
   or  u1 (OrCD_, C, D);
   or  u2 (OrAXB_, AX, B);
   not  u3 (AX, A);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO4AHS_D_F_Z_R,`AO4AHS_D_R_Z_F);
      (C -=> Z) = (`AO4AHS_C_F_Z_R,`AO4AHS_C_R_Z_F);
      (B -=> Z) = (`AO4AHS_B_F_Z_R,`AO4AHS_B_R_Z_F);
      (A +=> Z) = (`AO4AHS_A_R_Z_R,`AO4AHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO4AHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:06 and Version :1.1 //
 
//  START 
// CELL AO4AHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO4AHSP_D_F_Z_R 0.1
`define AO4AHSP_D_R_Z_F 0.1
`define AO4AHSP_C_F_Z_R 0.1
`define AO4AHSP_C_R_Z_F 0.1
`define AO4AHSP_B_F_Z_R 0.1
`define AO4AHSP_B_R_Z_F 0.1
`define AO4AHSP_A_F_Z_F 0.1
`define AO4AHSP_A_R_Z_R 0.1

module AO4AHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAXB_, OrCD_);
   or  u1 (OrCD_, C, D);
   or  u2 (OrAXB_, AX, B);
   not  u3 (AX, A);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO4AHSP_D_F_Z_R,`AO4AHSP_D_R_Z_F);
      (C -=> Z) = (`AO4AHSP_C_F_Z_R,`AO4AHSP_C_R_Z_F);
      (B -=> Z) = (`AO4AHSP_B_F_Z_R,`AO4AHSP_B_R_Z_F);
      (A +=> Z) = (`AO4AHSP_A_R_Z_R,`AO4AHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO4AHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:06 and Version :1.1 //
 
//  START 
// CELL AO4AHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO4AHSX4_D_F_Z_R 0.1
`define AO4AHSX4_D_R_Z_F 0.1
`define AO4AHSX4_C_F_Z_R 0.1
`define AO4AHSX4_C_R_Z_F 0.1
`define AO4AHSX4_B_F_Z_R 0.1
`define AO4AHSX4_B_R_Z_F 0.1
`define AO4AHSX4_A_F_Z_F 0.1
`define AO4AHSX4_A_R_Z_R 0.1

module AO4AHSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAXB_, OrCD_);
   or  u1 (OrCD_, C, D);
   or  u2 (OrAXB_, AX, B);
   not  u3 (AX, A);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO4AHSX4_D_F_Z_R,`AO4AHSX4_D_R_Z_F);
      (C -=> Z) = (`AO4AHSX4_C_F_Z_R,`AO4AHSX4_C_R_Z_F);
      (B -=> Z) = (`AO4AHSX4_B_F_Z_R,`AO4AHSX4_B_R_Z_F);
      (A +=> Z) = (`AO4AHSX4_A_R_Z_R,`AO4AHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO4AHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:06 and Version :1.1 //
 
//  START 
// CELL AO4AHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO4AHSX8_D_F_Z_R 0.1
`define AO4AHSX8_D_R_Z_F 0.1
`define AO4AHSX8_C_F_Z_R 0.1
`define AO4AHSX8_C_R_Z_F 0.1
`define AO4AHSX8_B_F_Z_R 0.1
`define AO4AHSX8_B_R_Z_F 0.1
`define AO4AHSX8_A_F_Z_F 0.1
`define AO4AHSX8_A_R_Z_R 0.1

module AO4AHSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAXB_, OrCD_);
   or  u1 (OrCD_, C, D);
   or  u2 (OrAXB_, AX, B);
   not  u3 (AX, A);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO4AHSX8_D_F_Z_R,`AO4AHSX8_D_R_Z_F);
      (C -=> Z) = (`AO4AHSX8_C_F_Z_R,`AO4AHSX8_C_R_Z_F);
      (B -=> Z) = (`AO4AHSX8_B_F_Z_R,`AO4AHSX8_B_R_Z_F);
      (A +=> Z) = (`AO4AHSX8_A_R_Z_R,`AO4AHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO4AHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:06 and Version :1.1 //
 
//  START 
// CELL F_AO4AHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO4AHSP_D_F_Z_R 0.1
`define F_AO4AHSP_D_R_Z_F 0.1
`define F_AO4AHSP_C_F_Z_R 0.1
`define F_AO4AHSP_C_R_Z_F 0.1
`define F_AO4AHSP_B_F_Z_R 0.1
`define F_AO4AHSP_B_R_Z_F 0.1
`define F_AO4AHSP_A_F_Z_F 0.1
`define F_AO4AHSP_A_R_Z_R 0.1

module F_AO4AHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, OrAXB_, OrCD_);
   or  u1 (OrCD_, C, D);
   or  u2 (OrAXB_, AX, B);
   not  u3 (AX, A);


`ifdef functional
`else
   specify

      (D -=> Z) = (`F_AO4AHSP_D_F_Z_R,`F_AO4AHSP_D_R_Z_F);
      (C -=> Z) = (`F_AO4AHSP_C_F_Z_R,`F_AO4AHSP_C_R_Z_F);
      (B -=> Z) = (`F_AO4AHSP_B_F_Z_R,`F_AO4AHSP_B_R_Z_F);
      (A +=> Z) = (`F_AO4AHSP_A_R_Z_R,`F_AO4AHSP_A_F_Z_F);

   endspecify
`endif


endmodule // F_AO4AHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:06 and Version :1.1 //
 
//  START 
// CELL AO4ANHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO4ANHS_D_F_Z_F 0.1
`define AO4ANHS_D_R_Z_R 0.1
`define AO4ANHS_C_F_Z_F 0.1
`define AO4ANHS_C_R_Z_R 0.1
`define AO4ANHS_B_F_Z_F 0.1
`define AO4ANHS_B_R_Z_R 0.1
`define AO4ANHS_A_F_Z_R 0.1
`define AO4ANHS_A_R_Z_F 0.1

module AO4ANHS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAXB_, OrCD_);
   or  u1 (OrCD_, C, D);
   or  u2 (OrAXB_, AX, B);
   not  u3 (AX, A);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO4ANHS_D_R_Z_R,`AO4ANHS_D_F_Z_F);
      (C +=> Z) = (`AO4ANHS_C_R_Z_R,`AO4ANHS_C_F_Z_F);
      (B +=> Z) = (`AO4ANHS_B_R_Z_R,`AO4ANHS_B_F_Z_F);
      (A -=> Z) = (`AO4ANHS_A_F_Z_R,`AO4ANHS_A_R_Z_F);

   endspecify
`endif


endmodule // AO4ANHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:06 and Version :1.1 //
 
//  START 
// CELL AO4ANHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO4ANHSP_D_F_Z_F 0.1
`define AO4ANHSP_D_R_Z_R 0.1
`define AO4ANHSP_C_F_Z_F 0.1
`define AO4ANHSP_C_R_Z_R 0.1
`define AO4ANHSP_B_F_Z_F 0.1
`define AO4ANHSP_B_R_Z_R 0.1
`define AO4ANHSP_A_F_Z_R 0.1
`define AO4ANHSP_A_R_Z_F 0.1

module AO4ANHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAXB_, OrCD_);
   or  u1 (OrCD_, C, D);
   or  u2 (OrAXB_, AX, B);
   not  u3 (AX, A);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO4ANHSP_D_R_Z_R,`AO4ANHSP_D_F_Z_F);
      (C +=> Z) = (`AO4ANHSP_C_R_Z_R,`AO4ANHSP_C_F_Z_F);
      (B +=> Z) = (`AO4ANHSP_B_R_Z_R,`AO4ANHSP_B_F_Z_F);
      (A -=> Z) = (`AO4ANHSP_A_F_Z_R,`AO4ANHSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO4ANHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:06 and Version :1.1 //
 
//  START 
// CELL AO4ANHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO4ANHSX4_D_F_Z_F 0.1
`define AO4ANHSX4_D_R_Z_R 0.1
`define AO4ANHSX4_C_F_Z_F 0.1
`define AO4ANHSX4_C_R_Z_R 0.1
`define AO4ANHSX4_B_F_Z_F 0.1
`define AO4ANHSX4_B_R_Z_R 0.1
`define AO4ANHSX4_A_F_Z_R 0.1
`define AO4ANHSX4_A_R_Z_F 0.1

module AO4ANHSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAXB_, OrCD_);
   or  u1 (OrCD_, C, D);
   or  u2 (OrAXB_, AX, B);
   not  u3 (AX, A);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO4ANHSX4_D_R_Z_R,`AO4ANHSX4_D_F_Z_F);
      (C +=> Z) = (`AO4ANHSX4_C_R_Z_R,`AO4ANHSX4_C_F_Z_F);
      (B +=> Z) = (`AO4ANHSX4_B_R_Z_R,`AO4ANHSX4_B_F_Z_F);
      (A -=> Z) = (`AO4ANHSX4_A_F_Z_R,`AO4ANHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO4ANHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:06 and Version :1.1 //
 
//  START 
// CELL AO4ANHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO4ANHSX8_D_F_Z_F 0.1
`define AO4ANHSX8_D_R_Z_R 0.1
`define AO4ANHSX8_C_F_Z_F 0.1
`define AO4ANHSX8_C_R_Z_R 0.1
`define AO4ANHSX8_B_F_Z_F 0.1
`define AO4ANHSX8_B_R_Z_R 0.1
`define AO4ANHSX8_A_F_Z_R 0.1
`define AO4ANHSX8_A_R_Z_F 0.1

module AO4ANHSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAXB_, OrCD_);
   or  u1 (OrCD_, C, D);
   or  u2 (OrAXB_, AX, B);
   not  u3 (AX, A);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO4ANHSX8_D_R_Z_R,`AO4ANHSX8_D_F_Z_F);
      (C +=> Z) = (`AO4ANHSX8_C_R_Z_R,`AO4ANHSX8_C_F_Z_F);
      (B +=> Z) = (`AO4ANHSX8_B_R_Z_R,`AO4ANHSX8_B_F_Z_F);
      (A -=> Z) = (`AO4ANHSX8_A_F_Z_R,`AO4ANHSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AO4ANHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:06 and Version :1.1 //
 
//  START 
// CELL AO4NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO4NHS_D_F_Z_F 0.1
`define AO4NHS_D_R_Z_R 0.1
`define AO4NHS_C_F_Z_F 0.1
`define AO4NHS_C_R_Z_R 0.1
`define AO4NHS_B_F_Z_F 0.1
`define AO4NHS_B_R_Z_R 0.1
`define AO4NHS_A_F_Z_F 0.1
`define AO4NHS_A_R_Z_R 0.1

module AO4NHS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAB_, OrCD_);
   or  u1 (OrCD_, C, D);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO4NHS_D_R_Z_R,`AO4NHS_D_F_Z_F);
      (C +=> Z) = (`AO4NHS_C_R_Z_R,`AO4NHS_C_F_Z_F);
      (B +=> Z) = (`AO4NHS_B_R_Z_R,`AO4NHS_B_F_Z_F);
      (A +=> Z) = (`AO4NHS_A_R_Z_R,`AO4NHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO4NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:09 and Version :1.1 //
 
//  START 
// CELL AO4NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO4NHSP_D_F_Z_F 0.1
`define AO4NHSP_D_R_Z_R 0.1
`define AO4NHSP_C_F_Z_F 0.1
`define AO4NHSP_C_R_Z_R 0.1
`define AO4NHSP_B_F_Z_F 0.1
`define AO4NHSP_B_R_Z_R 0.1
`define AO4NHSP_A_F_Z_F 0.1
`define AO4NHSP_A_R_Z_R 0.1

module AO4NHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAB_, OrCD_);
   or  u1 (OrCD_, C, D);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO4NHSP_D_R_Z_R,`AO4NHSP_D_F_Z_F);
      (C +=> Z) = (`AO4NHSP_C_R_Z_R,`AO4NHSP_C_F_Z_F);
      (B +=> Z) = (`AO4NHSP_B_R_Z_R,`AO4NHSP_B_F_Z_F);
      (A +=> Z) = (`AO4NHSP_A_R_Z_R,`AO4NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO4NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:09 and Version :1.1 //
 
//  START 
// CELL AO4NHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO4NHSX4_D_F_Z_F 0.1
`define AO4NHSX4_D_R_Z_R 0.1
`define AO4NHSX4_C_F_Z_F 0.1
`define AO4NHSX4_C_R_Z_R 0.1
`define AO4NHSX4_B_F_Z_F 0.1
`define AO4NHSX4_B_R_Z_R 0.1
`define AO4NHSX4_A_F_Z_F 0.1
`define AO4NHSX4_A_R_Z_R 0.1

module AO4NHSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAB_, OrCD_);
   or  u1 (OrCD_, C, D);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO4NHSX4_D_R_Z_R,`AO4NHSX4_D_F_Z_F);
      (C +=> Z) = (`AO4NHSX4_C_R_Z_R,`AO4NHSX4_C_F_Z_F);
      (B +=> Z) = (`AO4NHSX4_B_R_Z_R,`AO4NHSX4_B_F_Z_F);
      (A +=> Z) = (`AO4NHSX4_A_R_Z_R,`AO4NHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO4NHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:09 and Version :1.1 //
 
//  START 
// CELL AO4NHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO4NHSX8_D_F_Z_F 0.1
`define AO4NHSX8_D_R_Z_R 0.1
`define AO4NHSX8_C_F_Z_F 0.1
`define AO4NHSX8_C_R_Z_R 0.1
`define AO4NHSX8_B_F_Z_F 0.1
`define AO4NHSX8_B_R_Z_R 0.1
`define AO4NHSX8_A_F_Z_F 0.1
`define AO4NHSX8_A_R_Z_R 0.1

module AO4NHSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (Z, OrAB_, OrCD_);
   or  u1 (OrCD_, C, D);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO4NHSX8_D_R_Z_R,`AO4NHSX8_D_F_Z_F);
      (C +=> Z) = (`AO4NHSX8_C_R_Z_R,`AO4NHSX8_C_F_Z_F);
      (B +=> Z) = (`AO4NHSX8_B_R_Z_R,`AO4NHSX8_B_F_Z_F);
      (A +=> Z) = (`AO4NHSX8_A_R_Z_R,`AO4NHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO4NHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:09 and Version :1.1 //
 
//  START 
// CELL AO5HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO5HS_C_F_Z_R 0.1
`define AO5HS_C_R_Z_F 0.1
`define AO5HS_B_F_Z_R 0.1
`define AO5HS_B_R_Z_F 0.1
`define AO5HS_A_F_Z_R 0.1
`define AO5HS_A_R_Z_F 0.1

module AO5HS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (AndAB_, A, B);
   or  u1 (OrAndAB_C_, AndAB_, C);
   or  u2 (OrAB_, A, B);
   nand  u3 (Z, OrAndAB_C_, OrAB_);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO5HS_C_F_Z_R,`AO5HS_C_R_Z_F);
      (B -=> Z) = (`AO5HS_B_F_Z_R,`AO5HS_B_R_Z_F);
      (A -=> Z) = (`AO5HS_A_F_Z_R,`AO5HS_A_R_Z_F);

   endspecify
`endif


endmodule // AO5HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:16 and Version :1.1 //
 
//  START 
// CELL AO5HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO5HSP_C_F_Z_R 0.1
`define AO5HSP_C_R_Z_F 0.1
`define AO5HSP_B_F_Z_R 0.1
`define AO5HSP_B_R_Z_F 0.1
`define AO5HSP_A_F_Z_R 0.1
`define AO5HSP_A_R_Z_F 0.1

module AO5HSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (AndAB_, A, B);
   or  u1 (OrAndAB_C_, AndAB_, C);
   or  u2 (OrAB_, A, B);
   nand  u3 (Z, OrAndAB_C_, OrAB_);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO5HSP_C_F_Z_R,`AO5HSP_C_R_Z_F);
      (B -=> Z) = (`AO5HSP_B_F_Z_R,`AO5HSP_B_R_Z_F);
      (A -=> Z) = (`AO5HSP_A_F_Z_R,`AO5HSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO5HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:16 and Version :1.1 //
 
//  START 
// CELL AO5HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO5HSX4_C_F_Z_R 0.1
`define AO5HSX4_C_R_Z_F 0.1
`define AO5HSX4_B_F_Z_R 0.1
`define AO5HSX4_B_R_Z_F 0.1
`define AO5HSX4_A_F_Z_R 0.1
`define AO5HSX4_A_R_Z_F 0.1

module AO5HSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (AndAB_, A, B);
   or  u1 (OrAndAB_C_, AndAB_, C);
   or  u2 (OrAB_, A, B);
   nand  u3 (Z, OrAndAB_C_, OrAB_);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO5HSX4_C_F_Z_R,`AO5HSX4_C_R_Z_F);
      (B -=> Z) = (`AO5HSX4_B_F_Z_R,`AO5HSX4_B_R_Z_F);
      (A -=> Z) = (`AO5HSX4_A_F_Z_R,`AO5HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO5HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:16 and Version :1.1 //
 
//  START 
// CELL AO5HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO5HSX8_C_F_Z_R 0.1
`define AO5HSX8_C_R_Z_F 0.1
`define AO5HSX8_B_F_Z_R 0.1
`define AO5HSX8_B_R_Z_F 0.1
`define AO5HSX8_A_F_Z_R 0.1
`define AO5HSX8_A_R_Z_F 0.1

module AO5HSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (AndAB_, A, B);
   or  u1 (OrAndAB_C_, AndAB_, C);
   or  u2 (OrAB_, A, B);
   nand  u3 (Z, OrAndAB_C_, OrAB_);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO5HSX8_C_F_Z_R,`AO5HSX8_C_R_Z_F);
      (B -=> Z) = (`AO5HSX8_B_F_Z_R,`AO5HSX8_B_R_Z_F);
      (A -=> Z) = (`AO5HSX8_A_F_Z_R,`AO5HSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AO5HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:16 and Version :1.1 //
 
//  START 
// CELL AO5AHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO5AHS_C_F_Z_R 0.1
`define AO5AHS_C_R_Z_F 0.1
`define AO5AHS_B_F_Z_R 0.1
`define AO5AHS_B_R_Z_F 0.1
`define AO5AHS_A_F_Z_F 0.1
`define AO5AHS_A_R_Z_R 0.1

module AO5AHS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, OrAndAXB_C_, OrAXB_);
   or  u1 (OrAXB_, AX, B);
   or  u2 (OrAndAXB_C_, AndAXB_, C);
   and  u3 (AndAXB_, AX, B);
   not  u4 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO5AHS_C_F_Z_R,`AO5AHS_C_R_Z_F);
      (B -=> Z) = (`AO5AHS_B_F_Z_R,`AO5AHS_B_R_Z_F);
      (A +=> Z) = (`AO5AHS_A_R_Z_R,`AO5AHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO5AHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:19 and Version :1.1 //
 
//  START 
// CELL AO5AHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO5AHSP_C_F_Z_R 0.1
`define AO5AHSP_C_R_Z_F 0.1
`define AO5AHSP_B_F_Z_R 0.1
`define AO5AHSP_B_R_Z_F 0.1
`define AO5AHSP_A_F_Z_F 0.1
`define AO5AHSP_A_R_Z_R 0.1

module AO5AHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, OrAndAXB_C_, OrAXB_);
   or  u1 (OrAXB_, AX, B);
   or  u2 (OrAndAXB_C_, AndAXB_, C);
   and  u3 (AndAXB_, AX, B);
   not  u4 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO5AHSP_C_F_Z_R,`AO5AHSP_C_R_Z_F);
      (B -=> Z) = (`AO5AHSP_B_F_Z_R,`AO5AHSP_B_R_Z_F);
      (A +=> Z) = (`AO5AHSP_A_R_Z_R,`AO5AHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO5AHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:19 and Version :1.1 //
 
//  START 
// CELL AO5AHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO5AHSX4_C_F_Z_R 0.1
`define AO5AHSX4_C_R_Z_F 0.1
`define AO5AHSX4_B_F_Z_R 0.1
`define AO5AHSX4_B_R_Z_F 0.1
`define AO5AHSX4_A_F_Z_F 0.1
`define AO5AHSX4_A_R_Z_R 0.1

module AO5AHSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, OrAndAXB_C_, OrAXB_);
   or  u1 (OrAXB_, AX, B);
   or  u2 (OrAndAXB_C_, AndAXB_, C);
   and  u3 (AndAXB_, AX, B);
   not  u4 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO5AHSX4_C_F_Z_R,`AO5AHSX4_C_R_Z_F);
      (B -=> Z) = (`AO5AHSX4_B_F_Z_R,`AO5AHSX4_B_R_Z_F);
      (A +=> Z) = (`AO5AHSX4_A_R_Z_R,`AO5AHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO5AHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:19 and Version :1.1 //
 
//  START 
// CELL AO5AHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO5AHSX8_C_F_Z_R 0.1
`define AO5AHSX8_C_R_Z_F 0.1
`define AO5AHSX8_B_F_Z_R 0.1
`define AO5AHSX8_B_R_Z_F 0.1
`define AO5AHSX8_A_F_Z_F 0.1
`define AO5AHSX8_A_R_Z_R 0.1

module AO5AHSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, OrAndAXB_C_, OrAXB_);
   or  u1 (OrAXB_, AX, B);
   or  u2 (OrAndAXB_C_, AndAXB_, C);
   and  u3 (AndAXB_, AX, B);
   not  u4 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO5AHSX8_C_F_Z_R,`AO5AHSX8_C_R_Z_F);
      (B -=> Z) = (`AO5AHSX8_B_F_Z_R,`AO5AHSX8_B_R_Z_F);
      (A +=> Z) = (`AO5AHSX8_A_R_Z_R,`AO5AHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO5AHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:19 and Version :1.1 //
 
//  START 
// CELL AO5ANHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO5ANHS_C_F_Z_F 0.1
`define AO5ANHS_C_R_Z_R 0.1
`define AO5ANHS_B_F_Z_F 0.1
`define AO5ANHS_B_R_Z_R 0.1
`define AO5ANHS_A_F_Z_R 0.1
`define AO5ANHS_A_R_Z_F 0.1

module AO5ANHS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AndOrBC_AX_, AndBC_);
   and  u1 (AndBC_, B, C);
   and  u2 (AndOrBC_AX_, OrBC_, AX);
   not  u3 (AX, A);
   or  u4 (OrBC_, B, C);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO5ANHS_C_R_Z_R,`AO5ANHS_C_F_Z_F);
      (B +=> Z) = (`AO5ANHS_B_R_Z_R,`AO5ANHS_B_F_Z_F);
      (A -=> Z) = (`AO5ANHS_A_F_Z_R,`AO5ANHS_A_R_Z_F);

   endspecify
`endif


endmodule // AO5ANHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:19 and Version :1.1 //
 
//  START 
// CELL AO5ANHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO5ANHSP_C_F_Z_F 0.1
`define AO5ANHSP_C_R_Z_R 0.1
`define AO5ANHSP_B_F_Z_F 0.1
`define AO5ANHSP_B_R_Z_R 0.1
`define AO5ANHSP_A_F_Z_R 0.1
`define AO5ANHSP_A_R_Z_F 0.1

module AO5ANHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AndOrBC_AX_, AndBC_);
   and  u1 (AndBC_, B, C);
   and  u2 (AndOrBC_AX_, OrBC_, AX);
   not  u3 (AX, A);
   or  u4 (OrBC_, B, C);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO5ANHSP_C_R_Z_R,`AO5ANHSP_C_F_Z_F);
      (B +=> Z) = (`AO5ANHSP_B_R_Z_R,`AO5ANHSP_B_F_Z_F);
      (A -=> Z) = (`AO5ANHSP_A_F_Z_R,`AO5ANHSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO5ANHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:19 and Version :1.1 //
 
//  START 
// CELL AO5ANHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO5ANHSX4_C_F_Z_F 0.1
`define AO5ANHSX4_C_R_Z_R 0.1
`define AO5ANHSX4_B_F_Z_F 0.1
`define AO5ANHSX4_B_R_Z_R 0.1
`define AO5ANHSX4_A_F_Z_R 0.1
`define AO5ANHSX4_A_R_Z_F 0.1

module AO5ANHSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AndOrBC_AX_, AndBC_);
   and  u1 (AndBC_, B, C);
   and  u2 (AndOrBC_AX_, OrBC_, AX);
   not  u3 (AX, A);
   or  u4 (OrBC_, B, C);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO5ANHSX4_C_R_Z_R,`AO5ANHSX4_C_F_Z_F);
      (B +=> Z) = (`AO5ANHSX4_B_R_Z_R,`AO5ANHSX4_B_F_Z_F);
      (A -=> Z) = (`AO5ANHSX4_A_F_Z_R,`AO5ANHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO5ANHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:19 and Version :1.1 //
 
//  START 
// CELL AO5ANHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO5ANHSX8_C_F_Z_F 0.1
`define AO5ANHSX8_C_R_Z_R 0.1
`define AO5ANHSX8_B_F_Z_F 0.1
`define AO5ANHSX8_B_R_Z_R 0.1
`define AO5ANHSX8_A_F_Z_R 0.1
`define AO5ANHSX8_A_R_Z_F 0.1

module AO5ANHSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AndOrBC_AX_, AndBC_);
   and  u1 (AndBC_, B, C);
   and  u2 (AndOrBC_AX_, OrBC_, AX);
   not  u3 (AX, A);
   or  u4 (OrBC_, B, C);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO5ANHSX8_C_R_Z_R,`AO5ANHSX8_C_F_Z_F);
      (B +=> Z) = (`AO5ANHSX8_B_R_Z_R,`AO5ANHSX8_B_F_Z_F);
      (A -=> Z) = (`AO5ANHSX8_A_F_Z_R,`AO5ANHSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AO5ANHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:19 and Version :1.1 //
 
//  START 
// CELL AO5NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO5NHS_C_F_Z_F 0.1
`define AO5NHS_C_R_Z_R 0.1
`define AO5NHS_B_F_Z_F 0.1
`define AO5NHS_B_R_Z_R 0.1
`define AO5NHS_A_F_Z_F 0.1
`define AO5NHS_A_R_Z_R 0.1

module AO5NHS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AndOrBC_A_, AndBC_);
   and  u1 (AndBC_, B, C);
   and  u2 (AndOrBC_A_, OrBC_, A);
   or  u3 (OrBC_, B, C);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO5NHS_C_R_Z_R,`AO5NHS_C_F_Z_F);
      (B +=> Z) = (`AO5NHS_B_R_Z_R,`AO5NHS_B_F_Z_F);
      (A +=> Z) = (`AO5NHS_A_R_Z_R,`AO5NHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO5NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:21 and Version :1.1 //
 
//  START 
// CELL AO5NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO5NHSP_C_F_Z_F 0.1
`define AO5NHSP_C_R_Z_R 0.1
`define AO5NHSP_B_F_Z_F 0.1
`define AO5NHSP_B_R_Z_R 0.1
`define AO5NHSP_A_F_Z_F 0.1
`define AO5NHSP_A_R_Z_R 0.1

module AO5NHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AndOrBC_A_, AndBC_);
   and  u1 (AndBC_, B, C);
   and  u2 (AndOrBC_A_, OrBC_, A);
   or  u3 (OrBC_, B, C);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO5NHSP_C_R_Z_R,`AO5NHSP_C_F_Z_F);
      (B +=> Z) = (`AO5NHSP_B_R_Z_R,`AO5NHSP_B_F_Z_F);
      (A +=> Z) = (`AO5NHSP_A_R_Z_R,`AO5NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO5NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:21 and Version :1.1 //
 
//  START 
// CELL AO5NHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO5NHSX4_C_F_Z_F 0.1
`define AO5NHSX4_C_R_Z_R 0.1
`define AO5NHSX4_B_F_Z_F 0.1
`define AO5NHSX4_B_R_Z_R 0.1
`define AO5NHSX4_A_F_Z_F 0.1
`define AO5NHSX4_A_R_Z_R 0.1

module AO5NHSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AndOrBC_A_, AndBC_);
   and  u1 (AndBC_, B, C);
   and  u2 (AndOrBC_A_, OrBC_, A);
   or  u3 (OrBC_, B, C);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO5NHSX4_C_R_Z_R,`AO5NHSX4_C_F_Z_F);
      (B +=> Z) = (`AO5NHSX4_B_R_Z_R,`AO5NHSX4_B_F_Z_F);
      (A +=> Z) = (`AO5NHSX4_A_R_Z_R,`AO5NHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO5NHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:21 and Version :1.1 //
 
//  START 
// CELL AO5NHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO5NHSX8_C_F_Z_F 0.1
`define AO5NHSX8_C_R_Z_R 0.1
`define AO5NHSX8_B_F_Z_F 0.1
`define AO5NHSX8_B_R_Z_R 0.1
`define AO5NHSX8_A_F_Z_F 0.1
`define AO5NHSX8_A_R_Z_R 0.1

module AO5NHSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AndOrBC_A_, AndBC_);
   and  u1 (AndBC_, B, C);
   and  u2 (AndOrBC_A_, OrBC_, A);
   or  u3 (OrBC_, B, C);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO5NHSX8_C_R_Z_R,`AO5NHSX8_C_F_Z_F);
      (B +=> Z) = (`AO5NHSX8_B_R_Z_R,`AO5NHSX8_B_F_Z_F);
      (A +=> Z) = (`AO5NHSX8_A_R_Z_R,`AO5NHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO5NHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:21 and Version :1.1 //
 
//  START 
// CELL F_AO5NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO5NHSP_C_F_Z_F 0.1
`define F_AO5NHSP_C_R_Z_R 0.1
`define F_AO5NHSP_B_F_Z_F 0.1
`define F_AO5NHSP_B_R_Z_R 0.1
`define F_AO5NHSP_A_F_Z_F 0.1
`define F_AO5NHSP_A_R_Z_R 0.1

module F_AO5NHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AndOrBC_A_, AndBC_);
   and  u1 (AndBC_, B, C);
   and  u2 (AndOrBC_A_, OrBC_, A);
   or  u3 (OrBC_, B, C);


`ifdef functional
`else
   specify

      (C +=> Z) = (`F_AO5NHSP_C_R_Z_R,`F_AO5NHSP_C_F_Z_F);
      (B +=> Z) = (`F_AO5NHSP_B_R_Z_R,`F_AO5NHSP_B_F_Z_F);
      (A +=> Z) = (`F_AO5NHSP_A_R_Z_R,`F_AO5NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // F_AO5NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:21 and Version :1.1 //
 
//  START 
// CELL F_AO5NHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO5NHSX4_C_F_Z_F 0.1
`define F_AO5NHSX4_C_R_Z_R 0.1
`define F_AO5NHSX4_B_F_Z_F 0.1
`define F_AO5NHSX4_B_R_Z_R 0.1
`define F_AO5NHSX4_A_F_Z_F 0.1
`define F_AO5NHSX4_A_R_Z_R 0.1

module F_AO5NHSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AndOrBC_A_, AndBC_);
   and  u1 (AndBC_, B, C);
   and  u2 (AndOrBC_A_, OrBC_, A);
   or  u3 (OrBC_, B, C);


`ifdef functional
`else
   specify

      (C +=> Z) = (`F_AO5NHSX4_C_R_Z_R,`F_AO5NHSX4_C_F_Z_F);
      (B +=> Z) = (`F_AO5NHSX4_B_R_Z_R,`F_AO5NHSX4_B_F_Z_F);
      (A +=> Z) = (`F_AO5NHSX4_A_R_Z_R,`F_AO5NHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // F_AO5NHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:21 and Version :1.1 //
 
//  START 
// CELL AO6HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6HSX05_C_F_Z_R 0.1
`define AO6HSX05_C_R_Z_F 0.1
`define AO6HSX05_B_F_Z_R 0.1
`define AO6HSX05_B_R_Z_F 0.1
`define AO6HSX05_A_F_Z_R 0.1
`define AO6HSX05_A_R_Z_F 0.1

module AO6HSX05 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, AndAB_, C);
   and  u1 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO6HSX05_C_F_Z_R,`AO6HSX05_C_R_Z_F);
      (B -=> Z) = (`AO6HSX05_B_F_Z_R,`AO6HSX05_B_R_Z_F);
      (A -=> Z) = (`AO6HSX05_A_F_Z_R,`AO6HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // AO6HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:28 and Version :1.1 //
 
//  START 
// CELL AO6HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6HS_C_F_Z_R 0.1
`define AO6HS_C_R_Z_F 0.1
`define AO6HS_B_F_Z_R 0.1
`define AO6HS_B_R_Z_F 0.1
`define AO6HS_A_F_Z_R 0.1
`define AO6HS_A_R_Z_F 0.1

module AO6HS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, AndAB_, C);
   and  u1 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO6HS_C_F_Z_R,`AO6HS_C_R_Z_F);
      (B -=> Z) = (`AO6HS_B_F_Z_R,`AO6HS_B_R_Z_F);
      (A -=> Z) = (`AO6HS_A_F_Z_R,`AO6HS_A_R_Z_F);

   endspecify
`endif


endmodule // AO6HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:28 and Version :1.1 //
 
//  START 
// CELL AO6HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6HSP_C_F_Z_R 0.1
`define AO6HSP_C_R_Z_F 0.1
`define AO6HSP_B_F_Z_R 0.1
`define AO6HSP_B_R_Z_F 0.1
`define AO6HSP_A_F_Z_R 0.1
`define AO6HSP_A_R_Z_F 0.1

module AO6HSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, AndAB_, C);
   and  u1 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO6HSP_C_F_Z_R,`AO6HSP_C_R_Z_F);
      (B -=> Z) = (`AO6HSP_B_F_Z_R,`AO6HSP_B_R_Z_F);
      (A -=> Z) = (`AO6HSP_A_F_Z_R,`AO6HSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO6HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:28 and Version :1.1 //
 
//  START 
// CELL AO6HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6HSX4_C_F_Z_R 0.1
`define AO6HSX4_C_R_Z_F 0.1
`define AO6HSX4_B_F_Z_R 0.1
`define AO6HSX4_B_R_Z_F 0.1
`define AO6HSX4_A_F_Z_R 0.1
`define AO6HSX4_A_R_Z_F 0.1

module AO6HSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, AndAB_, C);
   and  u1 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO6HSX4_C_F_Z_R,`AO6HSX4_C_R_Z_F);
      (B -=> Z) = (`AO6HSX4_B_F_Z_R,`AO6HSX4_B_R_Z_F);
      (A -=> Z) = (`AO6HSX4_A_F_Z_R,`AO6HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO6HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:28 and Version :1.1 //
 
//  START 
// CELL AO6HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6HSX8_C_F_Z_R 0.1
`define AO6HSX8_C_R_Z_F 0.1
`define AO6HSX8_B_F_Z_R 0.1
`define AO6HSX8_B_R_Z_F 0.1
`define AO6HSX8_A_F_Z_R 0.1
`define AO6HSX8_A_R_Z_F 0.1

module AO6HSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, AndAB_, C);
   and  u1 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO6HSX8_C_F_Z_R,`AO6HSX8_C_R_Z_F);
      (B -=> Z) = (`AO6HSX8_B_F_Z_R,`AO6HSX8_B_R_Z_F);
      (A -=> Z) = (`AO6HSX8_A_F_Z_R,`AO6HSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AO6HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:28 and Version :1.1 //
 
//  START 
// CELL F_AO6HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO6HS_C_F_Z_R 0.1
`define F_AO6HS_C_R_Z_F 0.1
`define F_AO6HS_B_F_Z_R 0.1
`define F_AO6HS_B_R_Z_F 0.1
`define F_AO6HS_A_F_Z_R 0.1
`define F_AO6HS_A_R_Z_F 0.1

module F_AO6HS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, AndAB_, C);
   and  u1 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (C -=> Z) = (`F_AO6HS_C_F_Z_R,`F_AO6HS_C_R_Z_F);
      (B -=> Z) = (`F_AO6HS_B_F_Z_R,`F_AO6HS_B_R_Z_F);
      (A -=> Z) = (`F_AO6HS_A_F_Z_R,`F_AO6HS_A_R_Z_F);

   endspecify
`endif


endmodule // F_AO6HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:28 and Version :1.1 //
 
//  START 
// CELL F_AO6HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO6HSP_C_F_Z_R 0.1
`define F_AO6HSP_C_R_Z_F 0.1
`define F_AO6HSP_B_F_Z_R 0.1
`define F_AO6HSP_B_R_Z_F 0.1
`define F_AO6HSP_A_F_Z_R 0.1
`define F_AO6HSP_A_R_Z_F 0.1

module F_AO6HSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, AndAB_, C);
   and  u1 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (C -=> Z) = (`F_AO6HSP_C_F_Z_R,`F_AO6HSP_C_R_Z_F);
      (B -=> Z) = (`F_AO6HSP_B_F_Z_R,`F_AO6HSP_B_R_Z_F);
      (A -=> Z) = (`F_AO6HSP_A_F_Z_R,`F_AO6HSP_A_R_Z_F);

   endspecify
`endif


endmodule // F_AO6HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:28 and Version :1.1 //
 
//  START 
// CELL AO6AHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6AHS_C_F_Z_R 0.1
`define AO6AHS_C_R_Z_F 0.1
`define AO6AHS_B_F_Z_R 0.1
`define AO6AHS_B_R_Z_F 0.1
`define AO6AHS_A_F_Z_F 0.1
`define AO6AHS_A_R_Z_R 0.1

module AO6AHS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, AndAXB_, C);
   and  u1 (AndAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO6AHS_C_F_Z_R,`AO6AHS_C_R_Z_F);
      (B -=> Z) = (`AO6AHS_B_F_Z_R,`AO6AHS_B_R_Z_F);
      (A +=> Z) = (`AO6AHS_A_R_Z_R,`AO6AHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO6AHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:30 and Version :1.1 //
 
//  START 
// CELL AO6AHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6AHSP_C_F_Z_R 0.1
`define AO6AHSP_C_R_Z_F 0.1
`define AO6AHSP_B_F_Z_R 0.1
`define AO6AHSP_B_R_Z_F 0.1
`define AO6AHSP_A_F_Z_F 0.1
`define AO6AHSP_A_R_Z_R 0.1

module AO6AHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, AndAXB_, C);
   and  u1 (AndAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO6AHSP_C_F_Z_R,`AO6AHSP_C_R_Z_F);
      (B -=> Z) = (`AO6AHSP_B_F_Z_R,`AO6AHSP_B_R_Z_F);
      (A +=> Z) = (`AO6AHSP_A_R_Z_R,`AO6AHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO6AHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:30 and Version :1.1 //
 
//  START 
// CELL AO6AHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6AHSX4_C_F_Z_R 0.1
`define AO6AHSX4_C_R_Z_F 0.1
`define AO6AHSX4_B_F_Z_R 0.1
`define AO6AHSX4_B_R_Z_F 0.1
`define AO6AHSX4_A_F_Z_F 0.1
`define AO6AHSX4_A_R_Z_R 0.1

module AO6AHSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, AndAXB_, C);
   and  u1 (AndAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO6AHSX4_C_F_Z_R,`AO6AHSX4_C_R_Z_F);
      (B -=> Z) = (`AO6AHSX4_B_F_Z_R,`AO6AHSX4_B_R_Z_F);
      (A +=> Z) = (`AO6AHSX4_A_R_Z_R,`AO6AHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO6AHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:30 and Version :1.1 //
 
//  START 
// CELL AO6AHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6AHSX8_C_F_Z_R 0.1
`define AO6AHSX8_C_R_Z_F 0.1
`define AO6AHSX8_B_F_Z_R 0.1
`define AO6AHSX8_B_R_Z_F 0.1
`define AO6AHSX8_A_F_Z_F 0.1
`define AO6AHSX8_A_R_Z_R 0.1

module AO6AHSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, AndAXB_, C);
   and  u1 (AndAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO6AHSX8_C_F_Z_R,`AO6AHSX8_C_R_Z_F);
      (B -=> Z) = (`AO6AHSX8_B_F_Z_R,`AO6AHSX8_B_R_Z_F);
      (A +=> Z) = (`AO6AHSX8_A_R_Z_R,`AO6AHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO6AHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:30 and Version :1.1 //
 
//  START 
// CELL AO6ANHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6ANHS_C_F_Z_F 0.1
`define AO6ANHS_C_R_Z_R 0.1
`define AO6ANHS_B_F_Z_F 0.1
`define AO6ANHS_B_R_Z_R 0.1
`define AO6ANHS_A_F_Z_R 0.1
`define AO6ANHS_A_R_Z_F 0.1

module AO6ANHS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AndAXB_, C);
   and  u1 (AndAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO6ANHS_C_R_Z_R,`AO6ANHS_C_F_Z_F);
      (B +=> Z) = (`AO6ANHS_B_R_Z_R,`AO6ANHS_B_F_Z_F);
      (A -=> Z) = (`AO6ANHS_A_F_Z_R,`AO6ANHS_A_R_Z_F);

   endspecify
`endif


endmodule // AO6ANHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:30 and Version :1.1 //
 
//  START 
// CELL AO6ANHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6ANHSP_C_F_Z_F 0.1
`define AO6ANHSP_C_R_Z_R 0.1
`define AO6ANHSP_B_F_Z_F 0.1
`define AO6ANHSP_B_R_Z_R 0.1
`define AO6ANHSP_A_F_Z_R 0.1
`define AO6ANHSP_A_R_Z_F 0.1

module AO6ANHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AndAXB_, C);
   and  u1 (AndAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO6ANHSP_C_R_Z_R,`AO6ANHSP_C_F_Z_F);
      (B +=> Z) = (`AO6ANHSP_B_R_Z_R,`AO6ANHSP_B_F_Z_F);
      (A -=> Z) = (`AO6ANHSP_A_F_Z_R,`AO6ANHSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO6ANHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:30 and Version :1.1 //
 
//  START 
// CELL AO6ANHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6ANHSX4_C_F_Z_F 0.1
`define AO6ANHSX4_C_R_Z_R 0.1
`define AO6ANHSX4_B_F_Z_F 0.1
`define AO6ANHSX4_B_R_Z_R 0.1
`define AO6ANHSX4_A_F_Z_R 0.1
`define AO6ANHSX4_A_R_Z_F 0.1

module AO6ANHSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AndAXB_, C);
   and  u1 (AndAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO6ANHSX4_C_R_Z_R,`AO6ANHSX4_C_F_Z_F);
      (B +=> Z) = (`AO6ANHSX4_B_R_Z_R,`AO6ANHSX4_B_F_Z_F);
      (A -=> Z) = (`AO6ANHSX4_A_F_Z_R,`AO6ANHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO6ANHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:30 and Version :1.1 //
 
//  START 
// CELL AO6ANHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6ANHSX8_C_F_Z_F 0.1
`define AO6ANHSX8_C_R_Z_R 0.1
`define AO6ANHSX8_B_F_Z_F 0.1
`define AO6ANHSX8_B_R_Z_R 0.1
`define AO6ANHSX8_A_F_Z_R 0.1
`define AO6ANHSX8_A_R_Z_F 0.1

module AO6ANHSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AndAXB_, C);
   and  u1 (AndAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO6ANHSX8_C_R_Z_R,`AO6ANHSX8_C_F_Z_F);
      (B +=> Z) = (`AO6ANHSX8_B_R_Z_R,`AO6ANHSX8_B_F_Z_F);
      (A -=> Z) = (`AO6ANHSX8_A_F_Z_R,`AO6ANHSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AO6ANHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:30 and Version :1.1 //
 
//  START 
// CELL AO6CHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6CHS_C_F_Z_F 0.1
`define AO6CHS_C_R_Z_R 0.1
`define AO6CHS_B_F_Z_R 0.1
`define AO6CHS_B_R_Z_F 0.1
`define AO6CHS_A_F_Z_R 0.1
`define AO6CHS_A_R_Z_F 0.1

module AO6CHS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, AndAB_, CX);
   not  u1 (CX, C);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO6CHS_C_R_Z_R,`AO6CHS_C_F_Z_F);
      (B -=> Z) = (`AO6CHS_B_F_Z_R,`AO6CHS_B_R_Z_F);
      (A -=> Z) = (`AO6CHS_A_F_Z_R,`AO6CHS_A_R_Z_F);

   endspecify
`endif


endmodule // AO6CHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:37 and Version :1.1 //
 
//  START 
// CELL AO6CHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6CHSP_C_F_Z_F 0.1
`define AO6CHSP_C_R_Z_R 0.1
`define AO6CHSP_B_F_Z_R 0.1
`define AO6CHSP_B_R_Z_F 0.1
`define AO6CHSP_A_F_Z_R 0.1
`define AO6CHSP_A_R_Z_F 0.1

module AO6CHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, AndAB_, CX);
   not  u1 (CX, C);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO6CHSP_C_R_Z_R,`AO6CHSP_C_F_Z_F);
      (B -=> Z) = (`AO6CHSP_B_F_Z_R,`AO6CHSP_B_R_Z_F);
      (A -=> Z) = (`AO6CHSP_A_F_Z_R,`AO6CHSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO6CHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:37 and Version :1.1 //
 
//  START 
// CELL AO6CHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6CHSX4_C_F_Z_F 0.1
`define AO6CHSX4_C_R_Z_R 0.1
`define AO6CHSX4_B_F_Z_R 0.1
`define AO6CHSX4_B_R_Z_F 0.1
`define AO6CHSX4_A_F_Z_R 0.1
`define AO6CHSX4_A_R_Z_F 0.1

module AO6CHSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, AndAB_, CX);
   not  u1 (CX, C);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO6CHSX4_C_R_Z_R,`AO6CHSX4_C_F_Z_F);
      (B -=> Z) = (`AO6CHSX4_B_F_Z_R,`AO6CHSX4_B_R_Z_F);
      (A -=> Z) = (`AO6CHSX4_A_F_Z_R,`AO6CHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO6CHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:37 and Version :1.1 //
 
//  START 
// CELL AO6CHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6CHSX8_C_F_Z_F 0.1
`define AO6CHSX8_C_R_Z_R 0.1
`define AO6CHSX8_B_F_Z_R 0.1
`define AO6CHSX8_B_R_Z_F 0.1
`define AO6CHSX8_A_F_Z_R 0.1
`define AO6CHSX8_A_R_Z_F 0.1

module AO6CHSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, AndAB_, CX);
   not  u1 (CX, C);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO6CHSX8_C_R_Z_R,`AO6CHSX8_C_F_Z_F);
      (B -=> Z) = (`AO6CHSX8_B_F_Z_R,`AO6CHSX8_B_R_Z_F);
      (A -=> Z) = (`AO6CHSX8_A_F_Z_R,`AO6CHSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AO6CHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:37 and Version :1.1 //
 
//  START 
// CELL F_AO6CHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO6CHSP_C_F_Z_F 0.1
`define F_AO6CHSP_C_R_Z_R 0.1
`define F_AO6CHSP_B_F_Z_R 0.1
`define F_AO6CHSP_B_R_Z_F 0.1
`define F_AO6CHSP_A_F_Z_R 0.1
`define F_AO6CHSP_A_R_Z_F 0.1

module F_AO6CHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, AndAB_, CX);
   not  u1 (CX, C);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (C +=> Z) = (`F_AO6CHSP_C_R_Z_R,`F_AO6CHSP_C_F_Z_F);
      (B -=> Z) = (`F_AO6CHSP_B_F_Z_R,`F_AO6CHSP_B_R_Z_F);
      (A -=> Z) = (`F_AO6CHSP_A_F_Z_R,`F_AO6CHSP_A_R_Z_F);

   endspecify
`endif


endmodule // F_AO6CHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:37 and Version :1.1 //
 
//  START 
// CELL AO6CNHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6CNHS_C_F_Z_R 0.1
`define AO6CNHS_C_R_Z_F 0.1
`define AO6CNHS_B_F_Z_F 0.1
`define AO6CNHS_B_R_Z_R 0.1
`define AO6CNHS_A_F_Z_F 0.1
`define AO6CNHS_A_R_Z_R 0.1

module AO6CNHS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AndAB_, CX);
   not  u1 (CX, C);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO6CNHS_C_F_Z_R,`AO6CNHS_C_R_Z_F);
      (B +=> Z) = (`AO6CNHS_B_R_Z_R,`AO6CNHS_B_F_Z_F);
      (A +=> Z) = (`AO6CNHS_A_R_Z_R,`AO6CNHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO6CNHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:37 and Version :1.1 //
 
//  START 
// CELL AO6CNHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6CNHSP_C_F_Z_R 0.1
`define AO6CNHSP_C_R_Z_F 0.1
`define AO6CNHSP_B_F_Z_F 0.1
`define AO6CNHSP_B_R_Z_R 0.1
`define AO6CNHSP_A_F_Z_F 0.1
`define AO6CNHSP_A_R_Z_R 0.1

module AO6CNHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AndAB_, CX);
   not  u1 (CX, C);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO6CNHSP_C_F_Z_R,`AO6CNHSP_C_R_Z_F);
      (B +=> Z) = (`AO6CNHSP_B_R_Z_R,`AO6CNHSP_B_F_Z_F);
      (A +=> Z) = (`AO6CNHSP_A_R_Z_R,`AO6CNHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO6CNHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:37 and Version :1.1 //
 
//  START 
// CELL AO6CNHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6CNHSX4_C_F_Z_R 0.1
`define AO6CNHSX4_C_R_Z_F 0.1
`define AO6CNHSX4_B_F_Z_F 0.1
`define AO6CNHSX4_B_R_Z_R 0.1
`define AO6CNHSX4_A_F_Z_F 0.1
`define AO6CNHSX4_A_R_Z_R 0.1

module AO6CNHSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AndAB_, CX);
   not  u1 (CX, C);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO6CNHSX4_C_F_Z_R,`AO6CNHSX4_C_R_Z_F);
      (B +=> Z) = (`AO6CNHSX4_B_R_Z_R,`AO6CNHSX4_B_F_Z_F);
      (A +=> Z) = (`AO6CNHSX4_A_R_Z_R,`AO6CNHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO6CNHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:37 and Version :1.1 //
 
//  START 
// CELL AO6CNHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6CNHSX8_C_F_Z_R 0.1
`define AO6CNHSX8_C_R_Z_F 0.1
`define AO6CNHSX8_B_F_Z_F 0.1
`define AO6CNHSX8_B_R_Z_R 0.1
`define AO6CNHSX8_A_F_Z_F 0.1
`define AO6CNHSX8_A_R_Z_R 0.1

module AO6CNHSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AndAB_, CX);
   not  u1 (CX, C);
   and  u2 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO6CNHSX8_C_F_Z_R,`AO6CNHSX8_C_R_Z_F);
      (B +=> Z) = (`AO6CNHSX8_B_R_Z_R,`AO6CNHSX8_B_F_Z_F);
      (A +=> Z) = (`AO6CNHSX8_A_R_Z_R,`AO6CNHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO6CNHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:37 and Version :1.1 //
 
//  START 
// CELL AO6NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6NHS_C_F_Z_F 0.1
`define AO6NHS_C_R_Z_R 0.1
`define AO6NHS_B_F_Z_F 0.1
`define AO6NHS_B_R_Z_R 0.1
`define AO6NHS_A_F_Z_F 0.1
`define AO6NHS_A_R_Z_R 0.1

module AO6NHS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AndAB_, C);
   and  u1 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO6NHS_C_R_Z_R,`AO6NHS_C_F_Z_F);
      (B +=> Z) = (`AO6NHS_B_R_Z_R,`AO6NHS_B_F_Z_F);
      (A +=> Z) = (`AO6NHS_A_R_Z_R,`AO6NHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO6NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:39 and Version :1.1 //
 
//  START 
// CELL AO6NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6NHSP_C_F_Z_F 0.1
`define AO6NHSP_C_R_Z_R 0.1
`define AO6NHSP_B_F_Z_F 0.1
`define AO6NHSP_B_R_Z_R 0.1
`define AO6NHSP_A_F_Z_F 0.1
`define AO6NHSP_A_R_Z_R 0.1

module AO6NHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AndAB_, C);
   and  u1 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO6NHSP_C_R_Z_R,`AO6NHSP_C_F_Z_F);
      (B +=> Z) = (`AO6NHSP_B_R_Z_R,`AO6NHSP_B_F_Z_F);
      (A +=> Z) = (`AO6NHSP_A_R_Z_R,`AO6NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO6NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:39 and Version :1.1 //
 
//  START 
// CELL AO6NHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6NHSX4_C_F_Z_F 0.1
`define AO6NHSX4_C_R_Z_R 0.1
`define AO6NHSX4_B_F_Z_F 0.1
`define AO6NHSX4_B_R_Z_R 0.1
`define AO6NHSX4_A_F_Z_F 0.1
`define AO6NHSX4_A_R_Z_R 0.1

module AO6NHSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AndAB_, C);
   and  u1 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO6NHSX4_C_R_Z_R,`AO6NHSX4_C_F_Z_F);
      (B +=> Z) = (`AO6NHSX4_B_R_Z_R,`AO6NHSX4_B_F_Z_F);
      (A +=> Z) = (`AO6NHSX4_A_R_Z_R,`AO6NHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO6NHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:39 and Version :1.1 //
 
//  START 
// CELL AO6NHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO6NHSX8_C_F_Z_F 0.1
`define AO6NHSX8_C_R_Z_R 0.1
`define AO6NHSX8_B_F_Z_F 0.1
`define AO6NHSX8_B_R_Z_R 0.1
`define AO6NHSX8_A_F_Z_F 0.1
`define AO6NHSX8_A_R_Z_R 0.1

module AO6NHSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AndAB_, C);
   and  u1 (AndAB_, A, B);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO6NHSX8_C_R_Z_R,`AO6NHSX8_C_F_Z_F);
      (B +=> Z) = (`AO6NHSX8_B_R_Z_R,`AO6NHSX8_B_F_Z_F);
      (A +=> Z) = (`AO6NHSX8_A_R_Z_R,`AO6NHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO6NHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:39 and Version :1.1 //
 
//  START 
// CELL AO7HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7HSX05_C_F_Z_R 0.1
`define AO7HSX05_C_R_Z_F 0.1
`define AO7HSX05_B_F_Z_R 0.1
`define AO7HSX05_B_R_Z_F 0.1
`define AO7HSX05_A_F_Z_R 0.1
`define AO7HSX05_A_R_Z_F 0.1

module AO7HSX05 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, OrAB_, C);
   or  u1 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO7HSX05_C_F_Z_R,`AO7HSX05_C_R_Z_F);
      (B -=> Z) = (`AO7HSX05_B_F_Z_R,`AO7HSX05_B_R_Z_F);
      (A -=> Z) = (`AO7HSX05_A_F_Z_R,`AO7HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // AO7HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:46 and Version :1.1 //
 
//  START 
// CELL AO7HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7HS_C_F_Z_R 0.1
`define AO7HS_C_R_Z_F 0.1
`define AO7HS_B_F_Z_R 0.1
`define AO7HS_B_R_Z_F 0.1
`define AO7HS_A_F_Z_R 0.1
`define AO7HS_A_R_Z_F 0.1

module AO7HS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, OrAB_, C);
   or  u1 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO7HS_C_F_Z_R,`AO7HS_C_R_Z_F);
      (B -=> Z) = (`AO7HS_B_F_Z_R,`AO7HS_B_R_Z_F);
      (A -=> Z) = (`AO7HS_A_F_Z_R,`AO7HS_A_R_Z_F);

   endspecify
`endif


endmodule // AO7HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:46 and Version :1.1 //
 
//  START 
// CELL AO7HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7HSP_C_F_Z_R 0.1
`define AO7HSP_C_R_Z_F 0.1
`define AO7HSP_B_F_Z_R 0.1
`define AO7HSP_B_R_Z_F 0.1
`define AO7HSP_A_F_Z_R 0.1
`define AO7HSP_A_R_Z_F 0.1

module AO7HSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, OrAB_, C);
   or  u1 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO7HSP_C_F_Z_R,`AO7HSP_C_R_Z_F);
      (B -=> Z) = (`AO7HSP_B_F_Z_R,`AO7HSP_B_R_Z_F);
      (A -=> Z) = (`AO7HSP_A_F_Z_R,`AO7HSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO7HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:46 and Version :1.1 //
 
//  START 
// CELL AO7HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7HSX4_C_F_Z_R 0.1
`define AO7HSX4_C_R_Z_F 0.1
`define AO7HSX4_B_F_Z_R 0.1
`define AO7HSX4_B_R_Z_F 0.1
`define AO7HSX4_A_F_Z_R 0.1
`define AO7HSX4_A_R_Z_F 0.1

module AO7HSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, OrAB_, C);
   or  u1 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO7HSX4_C_F_Z_R,`AO7HSX4_C_R_Z_F);
      (B -=> Z) = (`AO7HSX4_B_F_Z_R,`AO7HSX4_B_R_Z_F);
      (A -=> Z) = (`AO7HSX4_A_F_Z_R,`AO7HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO7HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:46 and Version :1.1 //
 
//  START 
// CELL AO7HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7HSX8_C_F_Z_R 0.1
`define AO7HSX8_C_R_Z_F 0.1
`define AO7HSX8_B_F_Z_R 0.1
`define AO7HSX8_B_R_Z_F 0.1
`define AO7HSX8_A_F_Z_R 0.1
`define AO7HSX8_A_R_Z_F 0.1

module AO7HSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, OrAB_, C);
   or  u1 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO7HSX8_C_F_Z_R,`AO7HSX8_C_R_Z_F);
      (B -=> Z) = (`AO7HSX8_B_F_Z_R,`AO7HSX8_B_R_Z_F);
      (A -=> Z) = (`AO7HSX8_A_F_Z_R,`AO7HSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AO7HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:46 and Version :1.1 //
 
//  START 
// CELL F_AO7HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO7HS_C_F_Z_R 0.1
`define F_AO7HS_C_R_Z_F 0.1
`define F_AO7HS_B_F_Z_R 0.1
`define F_AO7HS_B_R_Z_F 0.1
`define F_AO7HS_A_F_Z_R 0.1
`define F_AO7HS_A_R_Z_F 0.1

module F_AO7HS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, OrAB_, C);
   or  u1 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (C -=> Z) = (`F_AO7HS_C_F_Z_R,`F_AO7HS_C_R_Z_F);
      (B -=> Z) = (`F_AO7HS_B_F_Z_R,`F_AO7HS_B_R_Z_F);
      (A -=> Z) = (`F_AO7HS_A_F_Z_R,`F_AO7HS_A_R_Z_F);

   endspecify
`endif


endmodule // F_AO7HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:46 and Version :1.1 //
 
//  START 
// CELL F_AO7HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO7HSP_C_F_Z_R 0.1
`define F_AO7HSP_C_R_Z_F 0.1
`define F_AO7HSP_B_F_Z_R 0.1
`define F_AO7HSP_B_R_Z_F 0.1
`define F_AO7HSP_A_F_Z_R 0.1
`define F_AO7HSP_A_R_Z_F 0.1

module F_AO7HSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, OrAB_, C);
   or  u1 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (C -=> Z) = (`F_AO7HSP_C_F_Z_R,`F_AO7HSP_C_R_Z_F);
      (B -=> Z) = (`F_AO7HSP_B_F_Z_R,`F_AO7HSP_B_R_Z_F);
      (A -=> Z) = (`F_AO7HSP_A_F_Z_R,`F_AO7HSP_A_R_Z_F);

   endspecify
`endif


endmodule // F_AO7HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:46 and Version :1.1 //
 
//  START 
// CELL AO7AHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7AHS_C_F_Z_R 0.1
`define AO7AHS_C_R_Z_F 0.1
`define AO7AHS_B_F_Z_R 0.1
`define AO7AHS_B_R_Z_F 0.1
`define AO7AHS_A_F_Z_F 0.1
`define AO7AHS_A_R_Z_R 0.1

module AO7AHS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, OrAXB_, C);
   or  u1 (OrAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO7AHS_C_F_Z_R,`AO7AHS_C_R_Z_F);
      (B -=> Z) = (`AO7AHS_B_F_Z_R,`AO7AHS_B_R_Z_F);
      (A +=> Z) = (`AO7AHS_A_R_Z_R,`AO7AHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO7AHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:49 and Version :1.1 //
 
//  START 
// CELL AO7AHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7AHSP_C_F_Z_R 0.1
`define AO7AHSP_C_R_Z_F 0.1
`define AO7AHSP_B_F_Z_R 0.1
`define AO7AHSP_B_R_Z_F 0.1
`define AO7AHSP_A_F_Z_F 0.1
`define AO7AHSP_A_R_Z_R 0.1

module AO7AHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, OrAXB_, C);
   or  u1 (OrAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO7AHSP_C_F_Z_R,`AO7AHSP_C_R_Z_F);
      (B -=> Z) = (`AO7AHSP_B_F_Z_R,`AO7AHSP_B_R_Z_F);
      (A +=> Z) = (`AO7AHSP_A_R_Z_R,`AO7AHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO7AHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:49 and Version :1.1 //
 
//  START 
// CELL AO7AHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7AHSX4_C_F_Z_R 0.1
`define AO7AHSX4_C_R_Z_F 0.1
`define AO7AHSX4_B_F_Z_R 0.1
`define AO7AHSX4_B_R_Z_F 0.1
`define AO7AHSX4_A_F_Z_F 0.1
`define AO7AHSX4_A_R_Z_R 0.1

module AO7AHSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, OrAXB_, C);
   or  u1 (OrAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO7AHSX4_C_F_Z_R,`AO7AHSX4_C_R_Z_F);
      (B -=> Z) = (`AO7AHSX4_B_F_Z_R,`AO7AHSX4_B_R_Z_F);
      (A +=> Z) = (`AO7AHSX4_A_R_Z_R,`AO7AHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO7AHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:49 and Version :1.1 //
 
//  START 
// CELL AO7AHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7AHSX8_C_F_Z_R 0.1
`define AO7AHSX8_C_R_Z_F 0.1
`define AO7AHSX8_B_F_Z_R 0.1
`define AO7AHSX8_B_R_Z_F 0.1
`define AO7AHSX8_A_F_Z_F 0.1
`define AO7AHSX8_A_R_Z_R 0.1

module AO7AHSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, OrAXB_, C);
   or  u1 (OrAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO7AHSX8_C_F_Z_R,`AO7AHSX8_C_R_Z_F);
      (B -=> Z) = (`AO7AHSX8_B_F_Z_R,`AO7AHSX8_B_R_Z_F);
      (A +=> Z) = (`AO7AHSX8_A_R_Z_R,`AO7AHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO7AHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:49 and Version :1.1 //
 
//  START 
// CELL F_AO7AHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO7AHSP_C_F_Z_R 0.1
`define F_AO7AHSP_C_R_Z_F 0.1
`define F_AO7AHSP_B_F_Z_R 0.1
`define F_AO7AHSP_B_R_Z_F 0.1
`define F_AO7AHSP_A_F_Z_F 0.1
`define F_AO7AHSP_A_R_Z_R 0.1

module F_AO7AHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, OrAXB_, C);
   or  u1 (OrAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`F_AO7AHSP_C_F_Z_R,`F_AO7AHSP_C_R_Z_F);
      (B -=> Z) = (`F_AO7AHSP_B_F_Z_R,`F_AO7AHSP_B_R_Z_F);
      (A +=> Z) = (`F_AO7AHSP_A_R_Z_R,`F_AO7AHSP_A_F_Z_F);

   endspecify
`endif


endmodule // F_AO7AHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:49 and Version :1.1 //
 
//  START 
// CELL AO7ANHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7ANHS_C_F_Z_F 0.1
`define AO7ANHS_C_R_Z_R 0.1
`define AO7ANHS_B_F_Z_F 0.1
`define AO7ANHS_B_R_Z_R 0.1
`define AO7ANHS_A_F_Z_R 0.1
`define AO7ANHS_A_R_Z_F 0.1

module AO7ANHS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (Z, OrAXB_, C);
   or  u1 (OrAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO7ANHS_C_R_Z_R,`AO7ANHS_C_F_Z_F);
      (B +=> Z) = (`AO7ANHS_B_R_Z_R,`AO7ANHS_B_F_Z_F);
      (A -=> Z) = (`AO7ANHS_A_F_Z_R,`AO7ANHS_A_R_Z_F);

   endspecify
`endif


endmodule // AO7ANHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:49 and Version :1.1 //
 
//  START 
// CELL AO7ANHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7ANHSP_C_F_Z_F 0.1
`define AO7ANHSP_C_R_Z_R 0.1
`define AO7ANHSP_B_F_Z_F 0.1
`define AO7ANHSP_B_R_Z_R 0.1
`define AO7ANHSP_A_F_Z_R 0.1
`define AO7ANHSP_A_R_Z_F 0.1

module AO7ANHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (Z, OrAXB_, C);
   or  u1 (OrAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO7ANHSP_C_R_Z_R,`AO7ANHSP_C_F_Z_F);
      (B +=> Z) = (`AO7ANHSP_B_R_Z_R,`AO7ANHSP_B_F_Z_F);
      (A -=> Z) = (`AO7ANHSP_A_F_Z_R,`AO7ANHSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO7ANHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:49 and Version :1.1 //
 
//  START 
// CELL AO7ANHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7ANHSX4_C_F_Z_F 0.1
`define AO7ANHSX4_C_R_Z_R 0.1
`define AO7ANHSX4_B_F_Z_F 0.1
`define AO7ANHSX4_B_R_Z_R 0.1
`define AO7ANHSX4_A_F_Z_R 0.1
`define AO7ANHSX4_A_R_Z_F 0.1

module AO7ANHSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (Z, OrAXB_, C);
   or  u1 (OrAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO7ANHSX4_C_R_Z_R,`AO7ANHSX4_C_F_Z_F);
      (B +=> Z) = (`AO7ANHSX4_B_R_Z_R,`AO7ANHSX4_B_F_Z_F);
      (A -=> Z) = (`AO7ANHSX4_A_F_Z_R,`AO7ANHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO7ANHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:49 and Version :1.1 //
 
//  START 
// CELL AO7ANHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7ANHSX8_C_F_Z_F 0.1
`define AO7ANHSX8_C_R_Z_R 0.1
`define AO7ANHSX8_B_F_Z_F 0.1
`define AO7ANHSX8_B_R_Z_R 0.1
`define AO7ANHSX8_A_F_Z_R 0.1
`define AO7ANHSX8_A_R_Z_F 0.1

module AO7ANHSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (Z, OrAXB_, C);
   or  u1 (OrAXB_, AX, B);
   not  u2 (AX, A);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO7ANHSX8_C_R_Z_R,`AO7ANHSX8_C_F_Z_F);
      (B +=> Z) = (`AO7ANHSX8_B_R_Z_R,`AO7ANHSX8_B_F_Z_F);
      (A -=> Z) = (`AO7ANHSX8_A_F_Z_R,`AO7ANHSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AO7ANHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:49 and Version :1.1 //
 
//  START 
// CELL AO7CHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7CHS_C_F_Z_F 0.1
`define AO7CHS_C_R_Z_R 0.1
`define AO7CHS_B_F_Z_R 0.1
`define AO7CHS_B_R_Z_F 0.1
`define AO7CHS_A_F_Z_R 0.1
`define AO7CHS_A_R_Z_F 0.1

module AO7CHS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, OrAB_, CX);
   not  u1 (CX, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO7CHS_C_R_Z_R,`AO7CHS_C_F_Z_F);
      (B -=> Z) = (`AO7CHS_B_F_Z_R,`AO7CHS_B_R_Z_F);
      (A -=> Z) = (`AO7CHS_A_F_Z_R,`AO7CHS_A_R_Z_F);

   endspecify
`endif


endmodule // AO7CHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:56 and Version :1.1 //
 
//  START 
// CELL AO7CHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7CHSP_C_F_Z_F 0.1
`define AO7CHSP_C_R_Z_R 0.1
`define AO7CHSP_B_F_Z_R 0.1
`define AO7CHSP_B_R_Z_F 0.1
`define AO7CHSP_A_F_Z_R 0.1
`define AO7CHSP_A_R_Z_F 0.1

module AO7CHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, OrAB_, CX);
   not  u1 (CX, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO7CHSP_C_R_Z_R,`AO7CHSP_C_F_Z_F);
      (B -=> Z) = (`AO7CHSP_B_F_Z_R,`AO7CHSP_B_R_Z_F);
      (A -=> Z) = (`AO7CHSP_A_F_Z_R,`AO7CHSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO7CHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:56 and Version :1.1 //
 
//  START 
// CELL AO7CHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7CHSX4_C_F_Z_F 0.1
`define AO7CHSX4_C_R_Z_R 0.1
`define AO7CHSX4_B_F_Z_R 0.1
`define AO7CHSX4_B_R_Z_F 0.1
`define AO7CHSX4_A_F_Z_R 0.1
`define AO7CHSX4_A_R_Z_F 0.1

module AO7CHSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, OrAB_, CX);
   not  u1 (CX, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO7CHSX4_C_R_Z_R,`AO7CHSX4_C_F_Z_F);
      (B -=> Z) = (`AO7CHSX4_B_F_Z_R,`AO7CHSX4_B_R_Z_F);
      (A -=> Z) = (`AO7CHSX4_A_F_Z_R,`AO7CHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO7CHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:56 and Version :1.1 //
 
//  START 
// CELL AO7CHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7CHSX8_C_F_Z_F 0.1
`define AO7CHSX8_C_R_Z_R 0.1
`define AO7CHSX8_B_F_Z_R 0.1
`define AO7CHSX8_B_R_Z_F 0.1
`define AO7CHSX8_A_F_Z_R 0.1
`define AO7CHSX8_A_R_Z_F 0.1

module AO7CHSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, OrAB_, CX);
   not  u1 (CX, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO7CHSX8_C_R_Z_R,`AO7CHSX8_C_F_Z_F);
      (B -=> Z) = (`AO7CHSX8_B_F_Z_R,`AO7CHSX8_B_R_Z_F);
      (A -=> Z) = (`AO7CHSX8_A_F_Z_R,`AO7CHSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AO7CHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:56 and Version :1.1 //
 
//  START 
// CELL F_AO7CHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO7CHS_C_F_Z_F 0.1
`define F_AO7CHS_C_R_Z_R 0.1
`define F_AO7CHS_B_F_Z_R 0.1
`define F_AO7CHS_B_R_Z_F 0.1
`define F_AO7CHS_A_F_Z_R 0.1
`define F_AO7CHS_A_R_Z_F 0.1

module F_AO7CHS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, OrAB_, CX);
   not  u1 (CX, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (C +=> Z) = (`F_AO7CHS_C_R_Z_R,`F_AO7CHS_C_F_Z_F);
      (B -=> Z) = (`F_AO7CHS_B_F_Z_R,`F_AO7CHS_B_R_Z_F);
      (A -=> Z) = (`F_AO7CHS_A_F_Z_R,`F_AO7CHS_A_R_Z_F);

   endspecify
`endif


endmodule // F_AO7CHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:56 and Version :1.1 //
 
//  START 
// CELL F_AO7CHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_AO7CHSP_C_F_Z_F 0.1
`define F_AO7CHSP_C_R_Z_R 0.1
`define F_AO7CHSP_B_F_Z_R 0.1
`define F_AO7CHSP_B_R_Z_F 0.1
`define F_AO7CHSP_A_F_Z_R 0.1
`define F_AO7CHSP_A_R_Z_F 0.1

module F_AO7CHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, OrAB_, CX);
   not  u1 (CX, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (C +=> Z) = (`F_AO7CHSP_C_R_Z_R,`F_AO7CHSP_C_F_Z_F);
      (B -=> Z) = (`F_AO7CHSP_B_F_Z_R,`F_AO7CHSP_B_R_Z_F);
      (A -=> Z) = (`F_AO7CHSP_A_F_Z_R,`F_AO7CHSP_A_R_Z_F);

   endspecify
`endif


endmodule // F_AO7CHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:56 and Version :1.1 //
 
//  START 
// CELL AO7CNHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7CNHS_C_F_Z_R 0.1
`define AO7CNHS_C_R_Z_F 0.1
`define AO7CNHS_B_F_Z_F 0.1
`define AO7CNHS_B_R_Z_R 0.1
`define AO7CNHS_A_F_Z_F 0.1
`define AO7CNHS_A_R_Z_R 0.1

module AO7CNHS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (Z, OrAB_, CX);
   not  u1 (CX, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO7CNHS_C_F_Z_R,`AO7CNHS_C_R_Z_F);
      (B +=> Z) = (`AO7CNHS_B_R_Z_R,`AO7CNHS_B_F_Z_F);
      (A +=> Z) = (`AO7CNHS_A_R_Z_R,`AO7CNHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO7CNHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:56 and Version :1.1 //
 
//  START 
// CELL AO7CNHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7CNHSP_C_F_Z_R 0.1
`define AO7CNHSP_C_R_Z_F 0.1
`define AO7CNHSP_B_F_Z_F 0.1
`define AO7CNHSP_B_R_Z_R 0.1
`define AO7CNHSP_A_F_Z_F 0.1
`define AO7CNHSP_A_R_Z_R 0.1

module AO7CNHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (Z, OrAB_, CX);
   not  u1 (CX, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO7CNHSP_C_F_Z_R,`AO7CNHSP_C_R_Z_F);
      (B +=> Z) = (`AO7CNHSP_B_R_Z_R,`AO7CNHSP_B_F_Z_F);
      (A +=> Z) = (`AO7CNHSP_A_R_Z_R,`AO7CNHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO7CNHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:56 and Version :1.1 //
 
//  START 
// CELL AO7CNHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7CNHSX4_C_F_Z_R 0.1
`define AO7CNHSX4_C_R_Z_F 0.1
`define AO7CNHSX4_B_F_Z_F 0.1
`define AO7CNHSX4_B_R_Z_R 0.1
`define AO7CNHSX4_A_F_Z_F 0.1
`define AO7CNHSX4_A_R_Z_R 0.1

module AO7CNHSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (Z, OrAB_, CX);
   not  u1 (CX, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO7CNHSX4_C_F_Z_R,`AO7CNHSX4_C_R_Z_F);
      (B +=> Z) = (`AO7CNHSX4_B_R_Z_R,`AO7CNHSX4_B_F_Z_F);
      (A +=> Z) = (`AO7CNHSX4_A_R_Z_R,`AO7CNHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO7CNHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:56 and Version :1.1 //
 
//  START 
// CELL AO7CNHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7CNHSX8_C_F_Z_R 0.1
`define AO7CNHSX8_C_R_Z_F 0.1
`define AO7CNHSX8_B_F_Z_F 0.1
`define AO7CNHSX8_B_R_Z_R 0.1
`define AO7CNHSX8_A_F_Z_F 0.1
`define AO7CNHSX8_A_R_Z_R 0.1

module AO7CNHSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (Z, OrAB_, CX);
   not  u1 (CX, C);
   or  u2 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (C -=> Z) = (`AO7CNHSX8_C_F_Z_R,`AO7CNHSX8_C_R_Z_F);
      (B +=> Z) = (`AO7CNHSX8_B_R_Z_R,`AO7CNHSX8_B_F_Z_F);
      (A +=> Z) = (`AO7CNHSX8_A_R_Z_R,`AO7CNHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO7CNHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:12:56 and Version :1.1 //
 
//  START 
// CELL AO7NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7NHS_C_F_Z_F 0.1
`define AO7NHS_C_R_Z_R 0.1
`define AO7NHS_B_F_Z_F 0.1
`define AO7NHS_B_R_Z_R 0.1
`define AO7NHS_A_F_Z_F 0.1
`define AO7NHS_A_R_Z_R 0.1

module AO7NHS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (Z, OrAB_, C);
   or  u1 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO7NHS_C_R_Z_R,`AO7NHS_C_F_Z_F);
      (B +=> Z) = (`AO7NHS_B_R_Z_R,`AO7NHS_B_F_Z_F);
      (A +=> Z) = (`AO7NHS_A_R_Z_R,`AO7NHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO7NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:00 and Version :1.1 //
 
//  START 
// CELL AO7NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7NHSP_C_F_Z_F 0.1
`define AO7NHSP_C_R_Z_R 0.1
`define AO7NHSP_B_F_Z_F 0.1
`define AO7NHSP_B_R_Z_R 0.1
`define AO7NHSP_A_F_Z_F 0.1
`define AO7NHSP_A_R_Z_R 0.1

module AO7NHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (Z, OrAB_, C);
   or  u1 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO7NHSP_C_R_Z_R,`AO7NHSP_C_F_Z_F);
      (B +=> Z) = (`AO7NHSP_B_R_Z_R,`AO7NHSP_B_F_Z_F);
      (A +=> Z) = (`AO7NHSP_A_R_Z_R,`AO7NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO7NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:00 and Version :1.1 //
 
//  START 
// CELL AO7NHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7NHSX4_C_F_Z_F 0.1
`define AO7NHSX4_C_R_Z_R 0.1
`define AO7NHSX4_B_F_Z_F 0.1
`define AO7NHSX4_B_R_Z_R 0.1
`define AO7NHSX4_A_F_Z_F 0.1
`define AO7NHSX4_A_R_Z_R 0.1

module AO7NHSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (Z, OrAB_, C);
   or  u1 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO7NHSX4_C_R_Z_R,`AO7NHSX4_C_F_Z_F);
      (B +=> Z) = (`AO7NHSX4_B_R_Z_R,`AO7NHSX4_B_F_Z_F);
      (A +=> Z) = (`AO7NHSX4_A_R_Z_R,`AO7NHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO7NHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:00 and Version :1.1 //
 
//  START 
// CELL AO7NHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO7NHSX8_C_F_Z_F 0.1
`define AO7NHSX8_C_R_Z_R 0.1
`define AO7NHSX8_B_F_Z_F 0.1
`define AO7NHSX8_B_R_Z_R 0.1
`define AO7NHSX8_A_F_Z_F 0.1
`define AO7NHSX8_A_R_Z_R 0.1

module AO7NHSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   and  u0 (Z, OrAB_, C);
   or  u1 (OrAB_, A, B);


`ifdef functional
`else
   specify

      (C +=> Z) = (`AO7NHSX8_C_R_Z_R,`AO7NHSX8_C_F_Z_F);
      (B +=> Z) = (`AO7NHSX8_B_R_Z_R,`AO7NHSX8_B_F_Z_F);
      (A +=> Z) = (`AO7NHSX8_A_R_Z_R,`AO7NHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO7NHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:00 and Version :1.1 //
 
//  START 
// CELL AO8HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO8HSX05_D_F_Z_R 0.1
`define AO8HSX05_D_R_Z_F 0.1
`define AO8HSX05_C_F_Z_R 0.1
`define AO8HSX05_C_R_Z_F 0.1
`define AO8HSX05_B_F_Z_R 0.1
`define AO8HSX05_B_R_Z_F 0.1
`define AO8HSX05_A_F_Z_R 0.1
`define AO8HSX05_A_R_Z_F 0.1

module AO8HSX05 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (AndABC_, A, B, C);
   nor  u1 (Z, AndABC_, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO8HSX05_D_F_Z_R,`AO8HSX05_D_R_Z_F);
      (C -=> Z) = (`AO8HSX05_C_F_Z_R,`AO8HSX05_C_R_Z_F);
      (B -=> Z) = (`AO8HSX05_B_F_Z_R,`AO8HSX05_B_R_Z_F);
      (A -=> Z) = (`AO8HSX05_A_F_Z_R,`AO8HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // AO8HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:18 and Version :1.1 //
 
//  START 
// CELL AO8HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO8HS_D_F_Z_R 0.1
`define AO8HS_D_R_Z_F 0.1
`define AO8HS_C_F_Z_R 0.1
`define AO8HS_C_R_Z_F 0.1
`define AO8HS_B_F_Z_R 0.1
`define AO8HS_B_R_Z_F 0.1
`define AO8HS_A_F_Z_R 0.1
`define AO8HS_A_R_Z_F 0.1

module AO8HS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (AndABC_, A, B, C);
   nor  u1 (Z, AndABC_, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO8HS_D_F_Z_R,`AO8HS_D_R_Z_F);
      (C -=> Z) = (`AO8HS_C_F_Z_R,`AO8HS_C_R_Z_F);
      (B -=> Z) = (`AO8HS_B_F_Z_R,`AO8HS_B_R_Z_F);
      (A -=> Z) = (`AO8HS_A_F_Z_R,`AO8HS_A_R_Z_F);

   endspecify
`endif


endmodule // AO8HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:18 and Version :1.1 //
 
//  START 
// CELL AO8HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO8HSP_D_F_Z_R 0.1
`define AO8HSP_D_R_Z_F 0.1
`define AO8HSP_C_F_Z_R 0.1
`define AO8HSP_C_R_Z_F 0.1
`define AO8HSP_B_F_Z_R 0.1
`define AO8HSP_B_R_Z_F 0.1
`define AO8HSP_A_F_Z_R 0.1
`define AO8HSP_A_R_Z_F 0.1

module AO8HSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (AndABC_, A, B, C);
   nor  u1 (Z, AndABC_, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO8HSP_D_F_Z_R,`AO8HSP_D_R_Z_F);
      (C -=> Z) = (`AO8HSP_C_F_Z_R,`AO8HSP_C_R_Z_F);
      (B -=> Z) = (`AO8HSP_B_F_Z_R,`AO8HSP_B_R_Z_F);
      (A -=> Z) = (`AO8HSP_A_F_Z_R,`AO8HSP_A_R_Z_F);

   endspecify
`endif


endmodule // AO8HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:18 and Version :1.1 //
 
//  START 
// CELL AO8HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO8HSX4_D_F_Z_R 0.1
`define AO8HSX4_D_R_Z_F 0.1
`define AO8HSX4_C_F_Z_R 0.1
`define AO8HSX4_C_R_Z_F 0.1
`define AO8HSX4_B_F_Z_R 0.1
`define AO8HSX4_B_R_Z_F 0.1
`define AO8HSX4_A_F_Z_R 0.1
`define AO8HSX4_A_R_Z_F 0.1

module AO8HSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (AndABC_, A, B, C);
   nor  u1 (Z, AndABC_, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO8HSX4_D_F_Z_R,`AO8HSX4_D_R_Z_F);
      (C -=> Z) = (`AO8HSX4_C_F_Z_R,`AO8HSX4_C_R_Z_F);
      (B -=> Z) = (`AO8HSX4_B_F_Z_R,`AO8HSX4_B_R_Z_F);
      (A -=> Z) = (`AO8HSX4_A_F_Z_R,`AO8HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO8HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:18 and Version :1.1 //
 
//  START 
// CELL AO8HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO8HSX8_D_F_Z_R 0.1
`define AO8HSX8_D_R_Z_F 0.1
`define AO8HSX8_C_F_Z_R 0.1
`define AO8HSX8_C_R_Z_F 0.1
`define AO8HSX8_B_F_Z_R 0.1
`define AO8HSX8_B_R_Z_F 0.1
`define AO8HSX8_A_F_Z_R 0.1
`define AO8HSX8_A_R_Z_F 0.1

module AO8HSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (AndABC_, A, B, C);
   nor  u1 (Z, AndABC_, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`AO8HSX8_D_F_Z_R,`AO8HSX8_D_R_Z_F);
      (C -=> Z) = (`AO8HSX8_C_F_Z_R,`AO8HSX8_C_R_Z_F);
      (B -=> Z) = (`AO8HSX8_B_F_Z_R,`AO8HSX8_B_R_Z_F);
      (A -=> Z) = (`AO8HSX8_A_F_Z_R,`AO8HSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AO8HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:18 and Version :1.1 //
 
//  START 
// CELL AO8NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO8NHS_D_F_Z_F 0.1
`define AO8NHS_D_R_Z_R 0.1
`define AO8NHS_C_F_Z_F 0.1
`define AO8NHS_C_R_Z_R 0.1
`define AO8NHS_B_F_Z_F 0.1
`define AO8NHS_B_R_Z_R 0.1
`define AO8NHS_A_F_Z_F 0.1
`define AO8NHS_A_R_Z_R 0.1

module AO8NHS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (AndABC_, A, B, C);
   or  u1 (Z, AndABC_, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO8NHS_D_R_Z_R,`AO8NHS_D_F_Z_F);
      (C +=> Z) = (`AO8NHS_C_R_Z_R,`AO8NHS_C_F_Z_F);
      (B +=> Z) = (`AO8NHS_B_R_Z_R,`AO8NHS_B_F_Z_F);
      (A +=> Z) = (`AO8NHS_A_R_Z_R,`AO8NHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO8NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:18 and Version :1.1 //
 
//  START 
// CELL AO8NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO8NHSP_D_F_Z_F 0.1
`define AO8NHSP_D_R_Z_R 0.1
`define AO8NHSP_C_F_Z_F 0.1
`define AO8NHSP_C_R_Z_R 0.1
`define AO8NHSP_B_F_Z_F 0.1
`define AO8NHSP_B_R_Z_R 0.1
`define AO8NHSP_A_F_Z_F 0.1
`define AO8NHSP_A_R_Z_R 0.1

module AO8NHSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (AndABC_, A, B, C);
   or  u1 (Z, AndABC_, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO8NHSP_D_R_Z_R,`AO8NHSP_D_F_Z_F);
      (C +=> Z) = (`AO8NHSP_C_R_Z_R,`AO8NHSP_C_F_Z_F);
      (B +=> Z) = (`AO8NHSP_B_R_Z_R,`AO8NHSP_B_F_Z_F);
      (A +=> Z) = (`AO8NHSP_A_R_Z_R,`AO8NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO8NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:18 and Version :1.1 //
 
//  START 
// CELL AO8NHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO8NHSX4_D_F_Z_F 0.1
`define AO8NHSX4_D_R_Z_R 0.1
`define AO8NHSX4_C_F_Z_F 0.1
`define AO8NHSX4_C_R_Z_R 0.1
`define AO8NHSX4_B_F_Z_F 0.1
`define AO8NHSX4_B_R_Z_R 0.1
`define AO8NHSX4_A_F_Z_F 0.1
`define AO8NHSX4_A_R_Z_R 0.1

module AO8NHSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (AndABC_, A, B, C);
   or  u1 (Z, AndABC_, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO8NHSX4_D_R_Z_R,`AO8NHSX4_D_F_Z_F);
      (C +=> Z) = (`AO8NHSX4_C_R_Z_R,`AO8NHSX4_C_F_Z_F);
      (B +=> Z) = (`AO8NHSX4_B_R_Z_R,`AO8NHSX4_B_F_Z_F);
      (A +=> Z) = (`AO8NHSX4_A_R_Z_R,`AO8NHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO8NHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:18 and Version :1.1 //
 
//  START 
// CELL AO8NHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO8NHSX8_D_F_Z_F 0.1
`define AO8NHSX8_D_R_Z_R 0.1
`define AO8NHSX8_C_F_Z_F 0.1
`define AO8NHSX8_C_R_Z_R 0.1
`define AO8NHSX8_B_F_Z_F 0.1
`define AO8NHSX8_B_R_Z_R 0.1
`define AO8NHSX8_A_F_Z_F 0.1
`define AO8NHSX8_A_R_Z_R 0.1

module AO8NHSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   and  u0 (AndABC_, A, B, C);
   or  u1 (Z, AndABC_, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`AO8NHSX8_D_R_Z_R,`AO8NHSX8_D_F_Z_F);
      (C +=> Z) = (`AO8NHSX8_C_R_Z_R,`AO8NHSX8_C_F_Z_F);
      (B +=> Z) = (`AO8NHSX8_B_R_Z_R,`AO8NHSX8_B_F_Z_F);
      (A +=> Z) = (`AO8NHSX8_A_R_Z_R,`AO8NHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO8NHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:18 and Version :1.1 //
 
//  START 
// CELL AO9HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO9HSX05_E_F_Z_R 0.1
`define AO9HSX05_E_R_Z_F 0.1
`define AO9HSX05_D_F_Z_R 0.1
`define AO9HSX05_D_R_Z_F 0.1
`define AO9HSX05_C_F_Z_R 0.1
`define AO9HSX05_C_R_Z_F 0.1
`define AO9HSX05_B_F_Z_R 0.1
`define AO9HSX05_B_R_Z_F 0.1
`define AO9HSX05_A_F_Z_R 0.1
`define AO9HSX05_A_R_Z_F 0.1

module AO9HSX05 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndABC_, A, B, C);
   and  u1 (AndDE_, D, E);
   nor  u2 (Z, AndABC_, AndDE_);


`ifdef functional
`else
   specify

      (E -=> Z) = (`AO9HSX05_E_F_Z_R,`AO9HSX05_E_R_Z_F);
      (D -=> Z) = (`AO9HSX05_D_F_Z_R,`AO9HSX05_D_R_Z_F);
      (C -=> Z) = (`AO9HSX05_C_F_Z_R,`AO9HSX05_C_R_Z_F);
      (B -=> Z) = (`AO9HSX05_B_F_Z_R,`AO9HSX05_B_R_Z_F);
      (A -=> Z) = (`AO9HSX05_A_F_Z_R,`AO9HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // AO9HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:37 and Version :1.1 //
 
//  START 
// CELL AO9HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO9HS_E_F_Z_R 0.1
`define AO9HS_E_R_Z_F 0.1
`define AO9HS_D_F_Z_R 0.1
`define AO9HS_D_R_Z_F 0.1
`define AO9HS_C_F_Z_R 0.1
`define AO9HS_C_R_Z_F 0.1
`define AO9HS_B_F_Z_R 0.1
`define AO9HS_B_R_Z_F 0.1
`define AO9HS_A_F_Z_R 0.1
`define AO9HS_A_R_Z_F 0.1

module AO9HS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndABC_, A, B, C);
   and  u1 (AndDE_, D, E);
   nor  u2 (Z, AndABC_, AndDE_);


`ifdef functional
`else
   specify

      (E -=> Z) = (`AO9HS_E_F_Z_R,`AO9HS_E_R_Z_F);
      (D -=> Z) = (`AO9HS_D_F_Z_R,`AO9HS_D_R_Z_F);
      (C -=> Z) = (`AO9HS_C_F_Z_R,`AO9HS_C_R_Z_F);
      (B -=> Z) = (`AO9HS_B_F_Z_R,`AO9HS_B_R_Z_F);
      (A -=> Z) = (`AO9HS_A_F_Z_R,`AO9HS_A_R_Z_F);

   endspecify
`endif


endmodule // AO9HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:37 and Version :1.1 //
 
//  START 
// CELL AO9HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO9HSX4_E_F_Z_R 0.1
`define AO9HSX4_E_R_Z_F 0.1
`define AO9HSX4_D_F_Z_R 0.1
`define AO9HSX4_D_R_Z_F 0.1
`define AO9HSX4_C_F_Z_R 0.1
`define AO9HSX4_C_R_Z_F 0.1
`define AO9HSX4_B_F_Z_R 0.1
`define AO9HSX4_B_R_Z_F 0.1
`define AO9HSX4_A_F_Z_R 0.1
`define AO9HSX4_A_R_Z_F 0.1

module AO9HSX4 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndABC_, A, B, C);
   and  u1 (AndDE_, D, E);
   nor  u2 (Z, AndABC_, AndDE_);


`ifdef functional
`else
   specify

      (E -=> Z) = (`AO9HSX4_E_F_Z_R,`AO9HSX4_E_R_Z_F);
      (D -=> Z) = (`AO9HSX4_D_F_Z_R,`AO9HSX4_D_R_Z_F);
      (C -=> Z) = (`AO9HSX4_C_F_Z_R,`AO9HSX4_C_R_Z_F);
      (B -=> Z) = (`AO9HSX4_B_F_Z_R,`AO9HSX4_B_R_Z_F);
      (A -=> Z) = (`AO9HSX4_A_F_Z_R,`AO9HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // AO9HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:37 and Version :1.1 //
 
//  START 
// CELL AO9HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO9HSX8_E_F_Z_R 0.1
`define AO9HSX8_E_R_Z_F 0.1
`define AO9HSX8_D_F_Z_R 0.1
`define AO9HSX8_D_R_Z_F 0.1
`define AO9HSX8_C_F_Z_R 0.1
`define AO9HSX8_C_R_Z_F 0.1
`define AO9HSX8_B_F_Z_R 0.1
`define AO9HSX8_B_R_Z_F 0.1
`define AO9HSX8_A_F_Z_R 0.1
`define AO9HSX8_A_R_Z_F 0.1

module AO9HSX8 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndABC_, A, B, C);
   and  u1 (AndDE_, D, E);
   nor  u2 (Z, AndABC_, AndDE_);


`ifdef functional
`else
   specify

      (E -=> Z) = (`AO9HSX8_E_F_Z_R,`AO9HSX8_E_R_Z_F);
      (D -=> Z) = (`AO9HSX8_D_F_Z_R,`AO9HSX8_D_R_Z_F);
      (C -=> Z) = (`AO9HSX8_C_F_Z_R,`AO9HSX8_C_R_Z_F);
      (B -=> Z) = (`AO9HSX8_B_F_Z_R,`AO9HSX8_B_R_Z_F);
      (A -=> Z) = (`AO9HSX8_A_F_Z_R,`AO9HSX8_A_R_Z_F);

   endspecify
`endif


endmodule // AO9HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:37 and Version :1.1 //
 
//  START 
// CELL AO9NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO9NHS_E_F_Z_F 0.1
`define AO9NHS_E_R_Z_R 0.1
`define AO9NHS_D_F_Z_F 0.1
`define AO9NHS_D_R_Z_R 0.1
`define AO9NHS_C_F_Z_F 0.1
`define AO9NHS_C_R_Z_R 0.1
`define AO9NHS_B_F_Z_F 0.1
`define AO9NHS_B_R_Z_R 0.1
`define AO9NHS_A_F_Z_F 0.1
`define AO9NHS_A_R_Z_R 0.1

module AO9NHS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndABC_, A, B, C);
   and  u1 (AndDE_, D, E);
   or  u2 (Z, AndABC_, AndDE_);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO9NHS_E_R_Z_R,`AO9NHS_E_F_Z_F);
      (D +=> Z) = (`AO9NHS_D_R_Z_R,`AO9NHS_D_F_Z_F);
      (C +=> Z) = (`AO9NHS_C_R_Z_R,`AO9NHS_C_F_Z_F);
      (B +=> Z) = (`AO9NHS_B_R_Z_R,`AO9NHS_B_F_Z_F);
      (A +=> Z) = (`AO9NHS_A_R_Z_R,`AO9NHS_A_F_Z_F);

   endspecify
`endif


endmodule // AO9NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:37 and Version :1.1 //
 
//  START 
// CELL AO9NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO9NHSP_E_F_Z_F 0.1
`define AO9NHSP_E_R_Z_R 0.1
`define AO9NHSP_D_F_Z_F 0.1
`define AO9NHSP_D_R_Z_R 0.1
`define AO9NHSP_C_F_Z_F 0.1
`define AO9NHSP_C_R_Z_R 0.1
`define AO9NHSP_B_F_Z_F 0.1
`define AO9NHSP_B_R_Z_R 0.1
`define AO9NHSP_A_F_Z_F 0.1
`define AO9NHSP_A_R_Z_R 0.1

module AO9NHSP (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndABC_, A, B, C);
   and  u1 (AndDE_, D, E);
   or  u2 (Z, AndABC_, AndDE_);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO9NHSP_E_R_Z_R,`AO9NHSP_E_F_Z_F);
      (D +=> Z) = (`AO9NHSP_D_R_Z_R,`AO9NHSP_D_F_Z_F);
      (C +=> Z) = (`AO9NHSP_C_R_Z_R,`AO9NHSP_C_F_Z_F);
      (B +=> Z) = (`AO9NHSP_B_R_Z_R,`AO9NHSP_B_F_Z_F);
      (A +=> Z) = (`AO9NHSP_A_R_Z_R,`AO9NHSP_A_F_Z_F);

   endspecify
`endif


endmodule // AO9NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:37 and Version :1.1 //
 
//  START 
// CELL AO9NHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO9NHSX4_E_F_Z_F 0.1
`define AO9NHSX4_E_R_Z_R 0.1
`define AO9NHSX4_D_F_Z_F 0.1
`define AO9NHSX4_D_R_Z_R 0.1
`define AO9NHSX4_C_F_Z_F 0.1
`define AO9NHSX4_C_R_Z_R 0.1
`define AO9NHSX4_B_F_Z_F 0.1
`define AO9NHSX4_B_R_Z_R 0.1
`define AO9NHSX4_A_F_Z_F 0.1
`define AO9NHSX4_A_R_Z_R 0.1

module AO9NHSX4 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndABC_, A, B, C);
   and  u1 (AndDE_, D, E);
   or  u2 (Z, AndABC_, AndDE_);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO9NHSX4_E_R_Z_R,`AO9NHSX4_E_F_Z_F);
      (D +=> Z) = (`AO9NHSX4_D_R_Z_R,`AO9NHSX4_D_F_Z_F);
      (C +=> Z) = (`AO9NHSX4_C_R_Z_R,`AO9NHSX4_C_F_Z_F);
      (B +=> Z) = (`AO9NHSX4_B_R_Z_R,`AO9NHSX4_B_F_Z_F);
      (A +=> Z) = (`AO9NHSX4_A_R_Z_R,`AO9NHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // AO9NHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:37 and Version :1.1 //
 
//  START 
// CELL AO9NHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AO9NHSX8_E_F_Z_F 0.1
`define AO9NHSX8_E_R_Z_R 0.1
`define AO9NHSX8_D_F_Z_F 0.1
`define AO9NHSX8_D_R_Z_R 0.1
`define AO9NHSX8_C_F_Z_F 0.1
`define AO9NHSX8_C_R_Z_R 0.1
`define AO9NHSX8_B_F_Z_F 0.1
`define AO9NHSX8_B_R_Z_R 0.1
`define AO9NHSX8_A_F_Z_F 0.1
`define AO9NHSX8_A_R_Z_R 0.1

module AO9NHSX8 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   and  u0 (AndABC_, A, B, C);
   and  u1 (AndDE_, D, E);
   or  u2 (Z, AndABC_, AndDE_);


`ifdef functional
`else
   specify

      (E +=> Z) = (`AO9NHSX8_E_R_Z_R,`AO9NHSX8_E_F_Z_F);
      (D +=> Z) = (`AO9NHSX8_D_R_Z_R,`AO9NHSX8_D_F_Z_F);
      (C +=> Z) = (`AO9NHSX8_C_R_Z_R,`AO9NHSX8_C_F_Z_F);
      (B +=> Z) = (`AO9NHSX8_B_R_Z_R,`AO9NHSX8_B_F_Z_F);
      (A +=> Z) = (`AO9NHSX8_A_R_Z_R,`AO9NHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // AO9NHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:37 and Version :1.1 //
 
//  START 
// CELL AS01HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AS01HS_CI_F_CO_F 0.1
`define AS01HS_CI_R_CO_R 0.1
`define AS01HS_B_F_CO_F 0.1
`define AS01HS_B_R_CO_R 0.1
`define AS01HS_B_F_CO_R 0.1
`define AS01HS_B_R_CO_F 0.1
`define AS01HS_A_F_CO_F 0.1
`define AS01HS_A_R_CO_R 0.1
`define AS01HS_ADD_F_CO_F 0.1
`define AS01HS_ADD_R_CO_R 0.1
`define AS01HS_ADD_F_CO_R 0.1
`define AS01HS_ADD_R_CO_F 0.1
`define AS01HS_CI_F_S_F 0.1
`define AS01HS_CI_R_S_R 0.1
`define AS01HS_CI_F_S_R 0.1
`define AS01HS_CI_R_S_F 0.1
`define AS01HS_B_F_S_F 0.1
`define AS01HS_B_R_S_R 0.1
`define AS01HS_B_F_S_R 0.1
`define AS01HS_B_R_S_F 0.1
`define AS01HS_A_F_S_F 0.1
`define AS01HS_A_R_S_R 0.1
`define AS01HS_A_F_S_R 0.1
`define AS01HS_A_R_S_F 0.1
`define AS01HS_ADD_F_S_F 0.1
`define AS01HS_ADD_R_S_R 0.1
`define AS01HS_ADD_F_S_R 0.1
`define AS01HS_ADD_R_S_F 0.1

module AS01HS (S, CO, A, B, CI, ADD);

   output S;
   output CO;
   input ADD;
   input A;
   input B;
   input CI;


   or  u0 (S, AndADDABCI_, AndADDXAXBCI_, AndADDXABXCI_, AndADDAXBXCI_, AndADDXABCIX_, AndADDAXBCIX_, AndADDABXCIX_, AndADDXAXBXCIX_);
   and  u1 (AndADDXAXBXCIX_, ADDX, AX, BX, CIX);
   and  u2 (AndADDABXCIX_, ADD, A, BX, CIX);
   and  u3 (AndADDAXBCIX_, ADD, AX, B, CIX);
   and  u4 (AndADDXABCIX_, ADDX, A, B, CIX);
   not  u5 (CIX, CI);
   and  u6 (AndADDAXBXCI_, ADD, AX, BX, CI);
   and  u7 (AndADDXABXCI_, ADDX, A, BX, CI);
   not  u8 (BX, B);
   and  u9 (AndADDXAXBCI_, ADDX, AX, B, CI);
   not  u10 (AX, A);
   not  u11 (ADDX, ADD);
   and  u12 (AndADDABCI_, ADD, A, B, CI);
   or  u13 (CO, AndADDBCI_, AndACI_, AndADDXBXCI_, AndADDAB_, AndADDXABX_);
   and  u14 (AndADDXABX_, ADDX, A, BX);
   and  u15 (AndADDAB_, ADD, A, B);
   and  u16 (AndADDXBXCI_, ADDX, BX, CI);
   and  u17 (AndACI_, A, CI);
   and  u18 (AndADDBCI_, ADD, B, CI);


`ifdef functional
`else
   specify

      (CI +=> CO) = (`AS01HS_CI_R_CO_R,`AS01HS_CI_F_CO_F);
      if (ADD && !A && CI || ADD && A && !CI) (B +=> CO) = (`AS01HS_B_R_CO_R,`AS01HS_B_F_CO_F);
      if (!ADD && !A && CI || !ADD && A && !CI) (B -=> CO) = (`AS01HS_B_F_CO_R,`AS01HS_B_R_CO_F);
      (A +=> CO) = (`AS01HS_A_R_CO_R,`AS01HS_A_F_CO_F);
      if (!A && B && CI || A && B && !CI) (ADD +=> CO) = (`AS01HS_ADD_R_CO_R,`AS01HS_ADD_F_CO_F);
      if (!A && !B && CI || A && !B && !CI) (ADD -=> CO) = (`AS01HS_ADD_F_CO_R,`AS01HS_ADD_R_CO_F);
      if (ADD && A && B || !ADD && !A && B || !ADD && A && !B || ADD && !A && !B) (CI +=> S) = (`AS01HS_CI_R_S_R,`AS01HS_CI_F_S_F);
      if (!ADD && A && B || ADD && !A && B || ADD && A && !B || !ADD && !A && !B) (CI -=> S) = (`AS01HS_CI_F_S_R,`AS01HS_CI_R_S_F);
      if (ADD && A && CI || !ADD && !A && CI || !ADD && A && !CI || ADD && !A && !CI) (B +=> S) = (`AS01HS_B_R_S_R,`AS01HS_B_F_S_F);
      if (!ADD && A && CI || ADD && !A && CI || ADD && A && !CI || !ADD && !A && !CI) (B -=> S) = (`AS01HS_B_F_S_R,`AS01HS_B_R_S_F);
      if (ADD && B && CI || !ADD && !B && CI || !ADD && B && !CI || ADD && !B && !CI) (A +=> S) = (`AS01HS_A_R_S_R,`AS01HS_A_F_S_F);
      if (!ADD && B && CI || ADD && !B && CI || ADD && B && !CI || !ADD && !B && !CI) (A -=> S) = (`AS01HS_A_F_S_R,`AS01HS_A_R_S_F);
      if (A && B && CI || !A && !B && CI || !A && B && !CI || A && !B && !CI) (ADD +=> S) = (`AS01HS_ADD_R_S_R,`AS01HS_ADD_F_S_F);
      if (!A && B && CI || A && !B && CI || A && B && !CI || !A && !B && !CI) (ADD -=> S) = (`AS01HS_ADD_F_S_R,`AS01HS_ADD_R_S_F);

   endspecify
`endif


endmodule // AS01HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:43 and Version :1.1 //
 
//  START 
// CELL AS01HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define AS01HSP_CI_F_CO_F 0.1
`define AS01HSP_CI_R_CO_R 0.1
`define AS01HSP_B_F_CO_F 0.1
`define AS01HSP_B_R_CO_R 0.1
`define AS01HSP_B_F_CO_R 0.1
`define AS01HSP_B_R_CO_F 0.1
`define AS01HSP_A_F_CO_F 0.1
`define AS01HSP_A_R_CO_R 0.1
`define AS01HSP_ADD_F_CO_F 0.1
`define AS01HSP_ADD_R_CO_R 0.1
`define AS01HSP_ADD_F_CO_R 0.1
`define AS01HSP_ADD_R_CO_F 0.1
`define AS01HSP_CI_F_S_F 0.1
`define AS01HSP_CI_R_S_R 0.1
`define AS01HSP_CI_F_S_R 0.1
`define AS01HSP_CI_R_S_F 0.1
`define AS01HSP_B_F_S_F 0.1
`define AS01HSP_B_R_S_R 0.1
`define AS01HSP_B_F_S_R 0.1
`define AS01HSP_B_R_S_F 0.1
`define AS01HSP_A_F_S_F 0.1
`define AS01HSP_A_R_S_R 0.1
`define AS01HSP_A_F_S_R 0.1
`define AS01HSP_A_R_S_F 0.1
`define AS01HSP_ADD_F_S_F 0.1
`define AS01HSP_ADD_R_S_R 0.1
`define AS01HSP_ADD_F_S_R 0.1
`define AS01HSP_ADD_R_S_F 0.1

module AS01HSP (S, CO, A, B, CI, ADD);

   output S;
   output CO;
   input ADD;
   input A;
   input B;
   input CI;


   or  u0 (S, AndADDABCI_, AndADDXAXBCI_, AndADDXABXCI_, AndADDAXBXCI_, AndADDXABCIX_, AndADDAXBCIX_, AndADDABXCIX_, AndADDXAXBXCIX_);
   and  u1 (AndADDXAXBXCIX_, ADDX, AX, BX, CIX);
   and  u2 (AndADDABXCIX_, ADD, A, BX, CIX);
   and  u3 (AndADDAXBCIX_, ADD, AX, B, CIX);
   and  u4 (AndADDXABCIX_, ADDX, A, B, CIX);
   not  u5 (CIX, CI);
   and  u6 (AndADDAXBXCI_, ADD, AX, BX, CI);
   and  u7 (AndADDXABXCI_, ADDX, A, BX, CI);
   not  u8 (BX, B);
   and  u9 (AndADDXAXBCI_, ADDX, AX, B, CI);
   not  u10 (AX, A);
   not  u11 (ADDX, ADD);
   and  u12 (AndADDABCI_, ADD, A, B, CI);
   or  u13 (CO, AndADDBCI_, AndACI_, AndADDXBXCI_, AndADDAB_, AndADDXABX_);
   and  u14 (AndADDXABX_, ADDX, A, BX);
   and  u15 (AndADDAB_, ADD, A, B);
   and  u16 (AndADDXBXCI_, ADDX, BX, CI);
   and  u17 (AndACI_, A, CI);
   and  u18 (AndADDBCI_, ADD, B, CI);


`ifdef functional
`else
   specify

      (CI +=> CO) = (`AS01HSP_CI_R_CO_R,`AS01HSP_CI_F_CO_F);
      if (ADD && !A && CI || ADD && A && !CI) (B +=> CO) = (`AS01HSP_B_R_CO_R,`AS01HSP_B_F_CO_F);
      if (!ADD && !A && CI || !ADD && A && !CI) (B -=> CO) = (`AS01HSP_B_F_CO_R,`AS01HSP_B_R_CO_F);
      (A +=> CO) = (`AS01HSP_A_R_CO_R,`AS01HSP_A_F_CO_F);
      if (!A && B && CI || A && B && !CI) (ADD +=> CO) = (`AS01HSP_ADD_R_CO_R,`AS01HSP_ADD_F_CO_F);
      if (!A && !B && CI || A && !B && !CI) (ADD -=> CO) = (`AS01HSP_ADD_F_CO_R,`AS01HSP_ADD_R_CO_F);
      if (ADD && A && B || !ADD && !A && B || !ADD && A && !B || ADD && !A && !B) (CI +=> S) = (`AS01HSP_CI_R_S_R,`AS01HSP_CI_F_S_F);
      if (!ADD && A && B || ADD && !A && B || ADD && A && !B || !ADD && !A && !B) (CI -=> S) = (`AS01HSP_CI_F_S_R,`AS01HSP_CI_R_S_F);
      if (ADD && A && CI || !ADD && !A && CI || !ADD && A && !CI || ADD && !A && !CI) (B +=> S) = (`AS01HSP_B_R_S_R,`AS01HSP_B_F_S_F);
      if (!ADD && A && CI || ADD && !A && CI || ADD && A && !CI || !ADD && !A && !CI) (B -=> S) = (`AS01HSP_B_F_S_R,`AS01HSP_B_R_S_F);
      if (ADD && B && CI || !ADD && !B && CI || !ADD && B && !CI || ADD && !B && !CI) (A +=> S) = (`AS01HSP_A_R_S_R,`AS01HSP_A_F_S_F);
      if (!ADD && B && CI || ADD && !B && CI || ADD && B && !CI || !ADD && !B && !CI) (A -=> S) = (`AS01HSP_A_F_S_R,`AS01HSP_A_R_S_F);
      if (A && B && CI || !A && !B && CI || !A && B && !CI || A && !B && !CI) (ADD +=> S) = (`AS01HSP_ADD_R_S_R,`AS01HSP_ADD_F_S_F);
      if (!A && B && CI || A && !B && CI || A && B && !CI || !A && !B && !CI) (ADD -=> S) = (`AS01HSP_ADD_F_S_R,`AS01HSP_ADD_R_S_F);

   endspecify
`endif


endmodule // AS01HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:13:43 and Version :1.1 //
 
//  START 
// Cell BFHS

`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define BFHS_A_R_Z_R 0.1
`define BFHS_A_F_Z_F 0.1

module BFHS (Z, A);

	output Z;
	input A;

	buf    U1 (Z, A) ;


`ifdef functional
`else

	specify

		(A +=> Z) = (`BFHS_A_R_Z_R,`BFHS_A_F_Z_F);


	endspecify

`endif

endmodule // BFHS

`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine

// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START
 
// Cell BFHSP

`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define BFHSP_A_R_Z_R 0.1
`define BFHSP_A_F_Z_F 0.1

module BFHSP (Z, A);

	output Z;
	input A;

	buf    U1 (Z, A) ;


`ifdef functional
`else

	specify

		(A +=> Z) = (`BFHSP_A_R_Z_R,`BFHSP_A_F_Z_F);


	endspecify

`endif

endmodule // BFHSP

`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine

// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START
 
// Cell BFHSX3

`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define BFHSX3_A_R_Z_R 0.1
`define BFHSX3_A_F_Z_F 0.1

module BFHSX3 (Z, A);

	output Z;
	input A;

	buf    U1 (Z, A) ;


`ifdef functional
`else

	specify

		(A +=> Z) = (`BFHSX3_A_R_Z_R,`BFHSX3_A_F_Z_F);


	endspecify

`endif

endmodule // BFHSX3

`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine

// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START
 
// Cell BFHSX4

`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define BFHSX4_A_R_Z_R 0.1
`define BFHSX4_A_F_Z_F 0.1

module BFHSX4 (Z, A);

	output Z;
	input A;

	buf    U1 (Z, A) ;


`ifdef functional
`else

	specify

		(A +=> Z) = (`BFHSX4_A_R_Z_R,`BFHSX4_A_F_Z_F);


	endspecify

`endif

endmodule // BFHSX4

`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine

// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START
 
// Cell BFHSX5

`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define BFHSX5_A_R_Z_R 0.1
`define BFHSX5_A_F_Z_F 0.1

module BFHSX5 (Z, A);

	output Z;
	input A;

	buf    U1 (Z, A) ;


`ifdef functional
`else

	specify

		(A +=> Z) = (`BFHSX5_A_R_Z_R,`BFHSX5_A_F_Z_F);


	endspecify

`endif

endmodule // BFHSX5

`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine

// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START
 
// Cell BFHSX8

`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define BFHSX8_A_R_Z_R 0.1
`define BFHSX8_A_F_Z_F 0.1

module BFHSX8 (Z, A);

	output Z;
	input A;

	buf    U1 (Z, A) ;


`ifdef functional
`else

	specify

		(A +=> Z) = (`BFHSX8_A_R_Z_R,`BFHSX8_A_F_Z_F);


	endspecify

`endif

endmodule // BFHSX8

`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine

// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START
 
// Cell BFHSX16

`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define BFHSX16_A_R_Z_R 0.1
`define BFHSX16_A_F_Z_F 0.1

module BFHSX16 (Z, A);

	output Z;
	input A;

	buf    U1 (Z, A) ;


`ifdef functional
`else

	specify

		(A +=> Z) = (`BFHSX16_A_R_Z_R,`BFHSX16_A_F_Z_F);


	endspecify

`endif

endmodule // BFHSX16

`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine

// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START
 
// Cell BFHSX32

`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define BFHSX32_A_R_Z_R 0.1
`define BFHSX32_A_F_Z_F 0.1

module BFHSX32 (Z, A);

	output Z;
	input A;

	buf    U1 (Z, A) ;


`ifdef functional
`else

	specify

		(A +=> Z) = (`BFHSX32_A_R_Z_R,`BFHSX32_A_F_Z_F);


	endspecify

`endif

endmodule // BFHSX32

`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine

// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START
 
// Cell CTBUFHSP

`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define CTBUFHSP_A_R_Z_R 0.1
`define CTBUFHSP_A_F_Z_F 0.1

module CTBUFHSP (Z, A);

	output Z;
	input A;

	buf    U1 (Z, A) ;


`ifdef functional
`else

	specify

		(A +=> Z) = (`CTBUFHSP_A_R_Z_R,`CTBUFHSP_A_F_Z_F);


	endspecify

`endif

endmodule // CTBUFHSP

`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine

// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START
 
// Cell CTBUFHSX4

`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define CTBUFHSX4_A_R_Z_R 0.1
`define CTBUFHSX4_A_F_Z_F 0.1

module CTBUFHSX4 (Z, A);

	output Z;
	input A;

	buf    U1 (Z, A) ;


`ifdef functional
`else

	specify

		(A +=> Z) = (`CTBUFHSX4_A_R_Z_R,`CTBUFHSX4_A_F_Z_F);


	endspecify

`endif

endmodule // CTBUFHSX4

`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine

// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START
 
// Cell CTBUFHSX8

`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define CTBUFHSX8_A_R_Z_R 0.1
`define CTBUFHSX8_A_F_Z_F 0.1

module CTBUFHSX8 (Z, A);

	output Z;
	input A;

	buf    U1 (Z, A) ;


`ifdef functional
`else

	specify

		(A +=> Z) = (`CTBUFHSX8_A_R_Z_R,`CTBUFHSX8_A_F_Z_F);


	endspecify

`endif

endmodule // CTBUFHSX8

`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine

// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START
 
// Cell CTBUFHSX16

`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define CTBUFHSX16_A_R_Z_R 0.1
`define CTBUFHSX16_A_F_Z_F 0.1

module CTBUFHSX16 (Z, A);

	output Z;
	input A;

	buf    U1 (Z, A) ;


`ifdef functional
`else

	specify

		(A +=> Z) = (`CTBUFHSX16_A_R_Z_R,`CTBUFHSX16_A_F_Z_F);


	endspecify

`endif

endmodule // CTBUFHSX16

`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine

// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START
 
// Cell CTBUFHSX32

`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define CTBUFHSX32_A_R_Z_R 0.1
`define CTBUFHSX32_A_F_Z_F 0.1

module CTBUFHSX32 (Z, A);

	output Z;
	input A;

	buf    U1 (Z, A) ;


`ifdef functional
`else

	specify

		(A +=> Z) = (`CTBUFHSX32_A_R_Z_R,`CTBUFHSX32_A_F_Z_F);


	endspecify

`endif

endmodule // CTBUFHSX32

`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine

// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START
 
// Cell DLY05HS

`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define DLY05HS_A_R_Z_R 0.1
`define DLY05HS_A_F_Z_F 0.1

module DLY05HS (Z, A);

	output Z;
	input A;

	buf    U1 (Z, A) ;


`ifdef functional
`else

	specify

		(A +=> Z) = (`DLY05HS_A_R_Z_R,`DLY05HS_A_F_Z_F);


	endspecify

`endif

endmodule // DLY05HS

`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine

// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START
 
// Cell DLY05HSP

`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define DLY05HSP_A_R_Z_R 0.1
`define DLY05HSP_A_F_Z_F 0.1

module DLY05HSP (Z, A);

	output Z;
	input A;

	buf    U1 (Z, A) ;


`ifdef functional
`else

	specify

		(A +=> Z) = (`DLY05HSP_A_R_Z_R,`DLY05HSP_A_F_Z_F);


	endspecify

`endif

endmodule // DLY05HSP

`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine

// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START
 
// Cell DLY1HSP

`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define DLY1HSP_A_R_Z_R 0.1
`define DLY1HSP_A_F_Z_F 0.1

module DLY1HSP (Z, A);

	output Z;
	input A;

	buf    U1 (Z, A) ;


`ifdef functional
`else

	specify

		(A +=> Z) = (`DLY1HSP_A_R_Z_R,`DLY1HSP_A_F_Z_F);


	endspecify

`endif

endmodule // DLY1HSP

`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine

// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START
 
// Cell DLY2HSP

`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define DLY2HSP_A_R_Z_R 0.1
`define DLY2HSP_A_F_Z_F 0.1

module DLY2HSP (Z, A);

	output Z;
	input A;

	buf    U1 (Z, A) ;


`ifdef functional
`else

	specify

		(A +=> Z) = (`DLY2HSP_A_R_Z_R,`DLY2HSP_A_F_Z_F);


	endspecify

`endif

endmodule // DLY2HSP

`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine

// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START
 
// Cell DLY4HSP

`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define DLY4HSP_A_R_Z_R 0.1
`define DLY4HSP_A_F_Z_F 0.1

module DLY4HSP (Z, A);

	output Z;
	input A;

	buf    U1 (Z, A) ;


`ifdef functional
`else

	specify

		(A +=> Z) = (`DLY4HSP_A_R_Z_R,`DLY4HSP_A_F_Z_F);


	endspecify

`endif

endmodule // DLY4HSP

`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine

// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START
 
// Cell F_BFHSX16

`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define F_BFHSX16_A_R_Z_R 0.1
`define F_BFHSX16_A_F_Z_F 0.1

module F_BFHSX16 (Z, A);

	output Z;
	input A;

	buf    U1 (Z, A) ;


`ifdef functional
`else

	specify

		(A +=> Z) = (`F_BFHSX16_A_R_Z_R,`F_BFHSX16_A_F_Z_F);


	endspecify

`endif

endmodule // F_BFHSX16

`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine

// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START
 
// Cell F_BFHSX8

`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define F_BFHSX8_A_R_Z_R 0.1
`define F_BFHSX8_A_F_Z_F 0.1

module F_BFHSX8 (Z, A);

	output Z;
	input A;

	buf    U1 (Z, A) ;


`ifdef functional
`else

	specify

		(A +=> Z) = (`F_BFHSX8_A_R_Z_R,`F_BFHSX8_A_F_Z_F);


	endspecify

`endif

endmodule // F_BFHSX8

`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine

// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START
 
// Cell M_BFHSP

`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define M_BFHSP_A_R_Z_R 0.1
`define M_BFHSP_A_F_Z_F 0.1

module M_BFHSP (Z, A);

	output Z;
	input A;

	buf    U1 (Z, A) ;


`ifdef functional
`else

	specify

		(A +=> Z) = (`M_BFHSP_A_R_Z_R,`M_BFHSP_A_F_Z_F);


	endspecify

`endif

endmodule // M_BFHSP

`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine

// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START
 
// CELL BK1HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

module BK1HS (A);
 
   inout A;
 
   not (weak0, weak1)  u0 (A, ZI);
   not                   u1 (ZI, A);
 
`ifdef functional
`else
   specify
 
   endspecify
`endif

endmodule // BK1HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:06 and Version :1.1 //
 
//  START 
// CELL BK1SHS
 
`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 
 
`define BK1SHS_TE_R_A_R 0.1
`define BK1SHS_TE_F_A_F 0.1
 
module BK1SHS (TE, A);
 
   input TE;
   inout A;
 
`ifdef TETRAMAX
 
   rnmos (A, TE, TE);
   not (weak0, weak1)  u0 (A, ZI);
   not                   u1 (ZI, A);
 
`else
 
   not (weak0, weak1)  u0 (A, ZI);
   nor                   u1 (ZI, TE, A);
 
`endif
 
`ifdef functional
`else
   specify
 
      (TE +=> A) = (`BK1SHS_TE_R_A_R,`BK1SHS_TE_F_A_F);
 
   endspecify
`endif
 
endmodule // BK1SHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
// CELL BTSHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define BTSHS_E_F_Z_HZ 0.1
`define BTSHS_E_R_Z_ZH 0.1
`define BTSHS_E_F_Z_LZ 0.1
`define BTSHS_E_R_Z_ZL 0.1
`define BTSHS_A_F_Z_F 0.1
`define BTSHS_A_R_Z_R 0.1

module BTSHS (Z, A, E);

   output Z;
   input A;
   input E;


   bufif1  u0 (Z, A, E);


`ifdef functional
`else
   specify

      (A +=> Z) = (`BTSHS_A_R_Z_R,`BTSHS_A_F_Z_F);
      (E => Z) = (`BTSHS_E_R_Z_ZH,`BTSHS_E_R_Z_ZL,`BTSHS_E_F_Z_LZ,`BTSHS_E_R_Z_ZH,`BTSHS_E_F_Z_HZ,`BTSHS_E_R_Z_ZL);

   endspecify
`endif


endmodule // BTSHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:13 and Version :1.1 //
 
//  START
// CELL BTSHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define BTSHSP_E_F_Z_HZ 0.1
`define BTSHSP_E_R_Z_ZH 0.1
`define BTSHSP_E_F_Z_LZ 0.1
`define BTSHSP_E_R_Z_ZL 0.1
`define BTSHSP_A_F_Z_F 0.1
`define BTSHSP_A_R_Z_R 0.1

module BTSHSP (Z, A, E);

   output Z;
   input A;
   input E;


   bufif1  u0 (Z, A, E);


`ifdef functional
`else
   specify

      (A +=> Z) = (`BTSHSP_A_R_Z_R,`BTSHSP_A_F_Z_F);
      (E => Z) = (`BTSHSP_E_R_Z_ZH,`BTSHSP_E_R_Z_ZL,`BTSHSP_E_F_Z_LZ,`BTSHSP_E_R_Z_ZH,`BTSHSP_E_F_Z_HZ,`BTSHSP_E_R_Z_ZL);

   endspecify
`endif


endmodule // BTSHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:13 and Version :1.1 //
 
//  START
// CELL BTSHSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define BTSHSX3_E_F_Z_HZ 0.1
`define BTSHSX3_E_R_Z_ZH 0.1
`define BTSHSX3_E_F_Z_LZ 0.1
`define BTSHSX3_E_R_Z_ZL 0.1
`define BTSHSX3_A_F_Z_F 0.1
`define BTSHSX3_A_R_Z_R 0.1

module BTSHSX3 (Z, A, E);

   output Z;
   input A;
   input E;


   bufif1  u0 (Z, A, E);


`ifdef functional
`else
   specify

      (A +=> Z) = (`BTSHSX3_A_R_Z_R,`BTSHSX3_A_F_Z_F);
      (E => Z) = (`BTSHSX3_E_R_Z_ZH,`BTSHSX3_E_R_Z_ZL,`BTSHSX3_E_F_Z_LZ,`BTSHSX3_E_R_Z_ZH,`BTSHSX3_E_F_Z_HZ,`BTSHSX3_E_R_Z_ZL);

   endspecify
`endif


endmodule // BTSHSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:13 and Version :1.1 //
 
//  START
// CELL BTSHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define BTSHSX4_E_F_Z_HZ 0.1
`define BTSHSX4_E_R_Z_ZH 0.1
`define BTSHSX4_E_F_Z_LZ 0.1
`define BTSHSX4_E_R_Z_ZL 0.1
`define BTSHSX4_A_F_Z_F 0.1
`define BTSHSX4_A_R_Z_R 0.1

module BTSHSX4 (Z, A, E);

   output Z;
   input A;
   input E;


   bufif1  u0 (Z, A, E);


`ifdef functional
`else
   specify

      (A +=> Z) = (`BTSHSX4_A_R_Z_R,`BTSHSX4_A_F_Z_F);
      (E => Z) = (`BTSHSX4_E_R_Z_ZH,`BTSHSX4_E_R_Z_ZL,`BTSHSX4_E_F_Z_LZ,`BTSHSX4_E_R_Z_ZH,`BTSHSX4_E_F_Z_HZ,`BTSHSX4_E_R_Z_ZL);

   endspecify
`endif


endmodule // BTSHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:13 and Version :1.1 //
 
//  START
// CELL BTSHSX5

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define BTSHSX5_E_F_Z_HZ 0.1
`define BTSHSX5_E_R_Z_ZH 0.1
`define BTSHSX5_E_F_Z_LZ 0.1
`define BTSHSX5_E_R_Z_ZL 0.1
`define BTSHSX5_A_F_Z_F 0.1
`define BTSHSX5_A_R_Z_R 0.1

module BTSHSX5 (Z, A, E);

   output Z;
   input A;
   input E;


   bufif1  u0 (Z, A, E);


`ifdef functional
`else
   specify

      (A +=> Z) = (`BTSHSX5_A_R_Z_R,`BTSHSX5_A_F_Z_F);
      (E => Z) = (`BTSHSX5_E_R_Z_ZH,`BTSHSX5_E_R_Z_ZL,`BTSHSX5_E_F_Z_LZ,`BTSHSX5_E_R_Z_ZH,`BTSHSX5_E_F_Z_HZ,`BTSHSX5_E_R_Z_ZL);

   endspecify
`endif


endmodule // BTSHSX5
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:13 and Version :1.1 //
 
//  START
// CELL BTSHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define BTSHSX8_E_F_Z_HZ 0.1
`define BTSHSX8_E_R_Z_ZH 0.1
`define BTSHSX8_E_F_Z_LZ 0.1
`define BTSHSX8_E_R_Z_ZL 0.1
`define BTSHSX8_A_F_Z_F 0.1
`define BTSHSX8_A_R_Z_R 0.1

module BTSHSX8 (Z, A, E);

   output Z;
   input A;
   input E;


   bufif1  u0 (Z, A, E);


`ifdef functional
`else
   specify

      (A +=> Z) = (`BTSHSX8_A_R_Z_R,`BTSHSX8_A_F_Z_F);
      (E => Z) = (`BTSHSX8_E_R_Z_ZH,`BTSHSX8_E_R_Z_ZL,`BTSHSX8_E_F_Z_LZ,`BTSHSX8_E_R_Z_ZH,`BTSHSX8_E_F_Z_HZ,`BTSHSX8_E_R_Z_ZL);

   endspecify
`endif


endmodule // BTSHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:13 and Version :1.1 //
 
//  START
// CELL BTSHSX16

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define BTSHSX16_E_F_Z_HZ 0.1
`define BTSHSX16_E_R_Z_ZH 0.1
`define BTSHSX16_E_F_Z_LZ 0.1
`define BTSHSX16_E_R_Z_ZL 0.1
`define BTSHSX16_A_F_Z_F 0.1
`define BTSHSX16_A_R_Z_R 0.1

module BTSHSX16 (Z, A, E);

   output Z;
   input A;
   input E;


   bufif1  u0 (Z, A, E);


`ifdef functional
`else
   specify

      (A +=> Z) = (`BTSHSX16_A_R_Z_R,`BTSHSX16_A_F_Z_F);
      (E => Z) = (`BTSHSX16_E_R_Z_ZH,`BTSHSX16_E_R_Z_ZL,`BTSHSX16_E_F_Z_LZ,`BTSHSX16_E_R_Z_ZH,`BTSHSX16_E_F_Z_HZ,`BTSHSX16_E_R_Z_ZL);

   endspecify
`endif


endmodule // BTSHSX16
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:13 and Version :1.1 //
 
//  START
// CELL BTSHSX32

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define BTSHSX32_E_F_Z_HZ 0.1
`define BTSHSX32_E_R_Z_ZH 0.1
`define BTSHSX32_E_F_Z_LZ 0.1
`define BTSHSX32_E_R_Z_ZL 0.1
`define BTSHSX32_A_F_Z_F 0.1
`define BTSHSX32_A_R_Z_R 0.1

module BTSHSX32 (Z, A, E);

   output Z;
   input A;
   input E;


   bufif1  u0 (Z, A, E);


`ifdef functional
`else
   specify

      (A +=> Z) = (`BTSHSX32_A_R_Z_R,`BTSHSX32_A_F_Z_F);
      (E => Z) = (`BTSHSX32_E_R_Z_ZH,`BTSHSX32_E_R_Z_ZL,`BTSHSX32_E_F_Z_LZ,`BTSHSX32_E_R_Z_ZH,`BTSHSX32_E_F_Z_HZ,`BTSHSX32_E_R_Z_ZL);

   endspecify
`endif


endmodule // BTSHSX32
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:13 and Version :1.1 //
 
//  START
// CELL BTSENHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define BTSENHS_EN_F_Z_ZH 0.1
`define BTSENHS_EN_R_Z_HZ 0.1
`define BTSENHS_EN_F_Z_ZL 0.1
`define BTSENHS_EN_R_Z_LZ 0.1
`define BTSENHS_A_F_Z_F 0.1
`define BTSENHS_A_R_Z_R 0.1

module BTSENHS (Z, A, EN);

   output Z;
   input A;
   input EN;


   bufif0  u0 (Z, A, EN);


`ifdef functional
`else
   specify

      (A +=> Z) = (`BTSENHS_A_R_Z_R,`BTSENHS_A_F_Z_F);
      (EN => Z) = (`BTSENHS_EN_F_Z_ZH,`BTSENHS_EN_F_Z_ZL,`BTSENHS_EN_R_Z_LZ,`BTSENHS_EN_F_Z_ZH,`BTSENHS_EN_R_Z_HZ,`BTSENHS_EN_F_Z_ZL);

   endspecify
`endif


endmodule // BTSENHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:13 and Version :1.1 //
 
//  START 
// CELL BTSENHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define BTSENHSP_EN_F_Z_ZH 0.1
`define BTSENHSP_EN_R_Z_HZ 0.1
`define BTSENHSP_EN_F_Z_ZL 0.1
`define BTSENHSP_EN_R_Z_LZ 0.1
`define BTSENHSP_A_F_Z_F 0.1
`define BTSENHSP_A_R_Z_R 0.1

module BTSENHSP (Z, A, EN);

   output Z;
   input A;
   input EN;


   bufif0  u0 (Z, A, EN);


`ifdef functional
`else
   specify

      (A +=> Z) = (`BTSENHSP_A_R_Z_R,`BTSENHSP_A_F_Z_F);
      (EN => Z) = (`BTSENHSP_EN_F_Z_ZH,`BTSENHSP_EN_F_Z_ZL,`BTSENHSP_EN_R_Z_LZ,`BTSENHSP_EN_F_Z_ZH,`BTSENHSP_EN_R_Z_HZ,`BTSENHSP_EN_F_Z_ZL);

   endspecify
`endif


endmodule // BTSENHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:13 and Version :1.1 //
 
//  START 
// CELL BTSENHSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define BTSENHSX3_EN_F_Z_ZH 0.1
`define BTSENHSX3_EN_R_Z_HZ 0.1
`define BTSENHSX3_EN_F_Z_ZL 0.1
`define BTSENHSX3_EN_R_Z_LZ 0.1
`define BTSENHSX3_A_F_Z_F 0.1
`define BTSENHSX3_A_R_Z_R 0.1

module BTSENHSX3 (Z, A, EN);

   output Z;
   input A;
   input EN;


   bufif0  u0 (Z, A, EN);


`ifdef functional
`else
   specify

      (A +=> Z) = (`BTSENHSX3_A_R_Z_R,`BTSENHSX3_A_F_Z_F);
      (EN => Z) = (`BTSENHSX3_EN_F_Z_ZH,`BTSENHSX3_EN_F_Z_ZL,`BTSENHSX3_EN_R_Z_LZ,`BTSENHSX3_EN_F_Z_ZH,`BTSENHSX3_EN_R_Z_HZ,`BTSENHSX3_EN_F_Z_ZL);

   endspecify
`endif


endmodule // BTSENHSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:13 and Version :1.1 //
 
//  START 
// CELL BTSENHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define BTSENHSX4_EN_F_Z_ZH 0.1
`define BTSENHSX4_EN_R_Z_HZ 0.1
`define BTSENHSX4_EN_F_Z_ZL 0.1
`define BTSENHSX4_EN_R_Z_LZ 0.1
`define BTSENHSX4_A_F_Z_F 0.1
`define BTSENHSX4_A_R_Z_R 0.1

module BTSENHSX4 (Z, A, EN);

   output Z;
   input A;
   input EN;


   bufif0  u0 (Z, A, EN);


`ifdef functional
`else
   specify

      (A +=> Z) = (`BTSENHSX4_A_R_Z_R,`BTSENHSX4_A_F_Z_F);
      (EN => Z) = (`BTSENHSX4_EN_F_Z_ZH,`BTSENHSX4_EN_F_Z_ZL,`BTSENHSX4_EN_R_Z_LZ,`BTSENHSX4_EN_F_Z_ZH,`BTSENHSX4_EN_R_Z_HZ,`BTSENHSX4_EN_F_Z_ZL);

   endspecify
`endif


endmodule // BTSENHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:13 and Version :1.1 //
 
//  START 
// CELL BTSENHSX5

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define BTSENHSX5_EN_F_Z_ZH 0.1
`define BTSENHSX5_EN_R_Z_HZ 0.1
`define BTSENHSX5_EN_F_Z_ZL 0.1
`define BTSENHSX5_EN_R_Z_LZ 0.1
`define BTSENHSX5_A_F_Z_F 0.1
`define BTSENHSX5_A_R_Z_R 0.1

module BTSENHSX5 (Z, A, EN);

   output Z;
   input A;
   input EN;


   bufif0  u0 (Z, A, EN);


`ifdef functional
`else
   specify

      (A +=> Z) = (`BTSENHSX5_A_R_Z_R,`BTSENHSX5_A_F_Z_F);
      (EN => Z) = (`BTSENHSX5_EN_F_Z_ZH,`BTSENHSX5_EN_F_Z_ZL,`BTSENHSX5_EN_R_Z_LZ,`BTSENHSX5_EN_F_Z_ZH,`BTSENHSX5_EN_R_Z_HZ,`BTSENHSX5_EN_F_Z_ZL);

   endspecify
`endif


endmodule // BTSENHSX5
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:13 and Version :1.1 //
 
//  START 
// CELL BTSENHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define BTSENHSX8_EN_F_Z_ZH 0.1
`define BTSENHSX8_EN_R_Z_HZ 0.1
`define BTSENHSX8_EN_F_Z_ZL 0.1
`define BTSENHSX8_EN_R_Z_LZ 0.1
`define BTSENHSX8_A_F_Z_F 0.1
`define BTSENHSX8_A_R_Z_R 0.1

module BTSENHSX8 (Z, A, EN);

   output Z;
   input A;
   input EN;


   bufif0  u0 (Z, A, EN);


`ifdef functional
`else
   specify

      (A +=> Z) = (`BTSENHSX8_A_R_Z_R,`BTSENHSX8_A_F_Z_F);
      (EN => Z) = (`BTSENHSX8_EN_F_Z_ZH,`BTSENHSX8_EN_F_Z_ZL,`BTSENHSX8_EN_R_Z_LZ,`BTSENHSX8_EN_F_Z_ZH,`BTSENHSX8_EN_R_Z_HZ,`BTSENHSX8_EN_F_Z_ZL);

   endspecify
`endif


endmodule // BTSENHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:13 and Version :1.1 //
 
//  START 
// CELL BTSENHSX16

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define BTSENHSX16_EN_F_Z_ZH 0.1
`define BTSENHSX16_EN_R_Z_HZ 0.1
`define BTSENHSX16_EN_F_Z_ZL 0.1
`define BTSENHSX16_EN_R_Z_LZ 0.1
`define BTSENHSX16_A_F_Z_F 0.1
`define BTSENHSX16_A_R_Z_R 0.1

module BTSENHSX16 (Z, A, EN);

   output Z;
   input A;
   input EN;


   bufif0  u0 (Z, A, EN);


`ifdef functional
`else
   specify

      (A +=> Z) = (`BTSENHSX16_A_R_Z_R,`BTSENHSX16_A_F_Z_F);
      (EN => Z) = (`BTSENHSX16_EN_F_Z_ZH,`BTSENHSX16_EN_F_Z_ZL,`BTSENHSX16_EN_R_Z_LZ,`BTSENHSX16_EN_F_Z_ZH,`BTSENHSX16_EN_R_Z_HZ,`BTSENHSX16_EN_F_Z_ZL);

   endspecify
`endif


endmodule // BTSENHSX16
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:13 and Version :1.1 //
 
//  START 
// CELL BTSENHSX32

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define BTSENHSX32_EN_F_Z_ZH 0.1
`define BTSENHSX32_EN_R_Z_HZ 0.1
`define BTSENHSX32_EN_F_Z_ZL 0.1
`define BTSENHSX32_EN_R_Z_LZ 0.1
`define BTSENHSX32_A_F_Z_F 0.1
`define BTSENHSX32_A_R_Z_R 0.1

module BTSENHSX32 (Z, A, EN);

   output Z;
   input A;
   input EN;


   bufif0  u0 (Z, A, EN);


`ifdef functional
`else
   specify

      (A +=> Z) = (`BTSENHSX32_A_R_Z_R,`BTSENHSX32_A_F_Z_F);
      (EN => Z) = (`BTSENHSX32_EN_F_Z_ZH,`BTSENHSX32_EN_F_Z_ZL,`BTSENHSX32_EN_R_Z_LZ,`BTSENHSX32_EN_F_Z_ZH,`BTSENHSX32_EN_R_Z_HZ,`BTSENHSX32_EN_F_Z_ZL);

   endspecify
`endif


endmodule // BTSENHSX32
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:13 and Version :1.1 //
 
//  START 
// CELL CBUFLHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define CBUFLHS_CP_F_G_F 0.1
`define CBUFLHS_CP_R_G_R 0.1
`define CBUFLHS_E_CP_HOLD 0.1
`define CBUFLHS_E_CP_SETUP 0.1
`define CBUFLHS_TE_CP_HOLD 0.1
`define CBUFLHS_TE_CP_SETUP 0.1
`define CBUFLHS_CP_PWL 0.1


module CBUFLHS (G, CP, E, TE );

	output G;
	input CP;
	input E;
	input TE;

   reg NOTIFIER;

	or    u0 (INTERNAL1, E, TE) ;
	U_LD_N_NOTI u1 (IQ, INTERNAL1, CP , NOTIFIER) ;
	and    u2 (INTERNAL2, IQ, CP) ;
	buf    u3 (G, INTERNAL2) ;


`ifdef functional
`else
   not  (TEX, TE);
   not  (EX, E);

	specify

		(CP +=> G) = (`CBUFLHS_CP_R_G_R,`CBUFLHS_CP_F_G_F);
      $setuphold(posedge CP &&& EX , posedge TE, `CBUFLHS_TE_CP_SETUP, `CBUFLHS_TE_CP_HOLD, NOTIFIER);
      $setuphold(posedge CP &&& EX , negedge TE, `CBUFLHS_TE_CP_SETUP, `CBUFLHS_TE_CP_HOLD, NOTIFIER);
      $setuphold(posedge CP &&& TEX , posedge E, `CBUFLHS_E_CP_SETUP, `CBUFLHS_E_CP_HOLD, NOTIFIER);
      $setuphold(posedge CP &&& TEX , negedge E, `CBUFLHS_E_CP_SETUP, `CBUFLHS_E_CP_HOLD, NOTIFIER);
      $width(negedge CP, `CBUFLHS_CP_PWL, 0, NOTIFIER);


	endspecify

`endif

endmodule // CBUFLHS

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
 
//  START
// CELL CBUFLHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define CBUFLHSP_CP_F_G_F 0.1
`define CBUFLHSP_CP_R_G_R 0.1
`define CBUFLHSP_E_CP_HOLD 0.1
`define CBUFLHSP_E_CP_SETUP 0.1
`define CBUFLHSP_TE_CP_HOLD 0.1
`define CBUFLHSP_TE_CP_SETUP 0.1
`define CBUFLHSP_CP_PWL 0.1


module CBUFLHSP (G, CP, E, TE );

	output G;
	input CP;
	input E;
	input TE;

   reg NOTIFIER;

	or    u0 (INTERNAL1, E, TE) ;
	U_LD_N_NOTI u1 (IQ, INTERNAL1, CP , NOTIFIER) ;
	and    u2 (INTERNAL2, IQ, CP) ;
	buf    u3 (G, INTERNAL2) ;


`ifdef functional
`else
   not  (TEX, TE);
   not  (EX, E);

	specify

		(CP +=> G) = (`CBUFLHSP_CP_R_G_R,`CBUFLHSP_CP_F_G_F);
      $setuphold(posedge CP &&& EX , posedge TE, `CBUFLHSP_TE_CP_SETUP, `CBUFLHSP_TE_CP_HOLD, NOTIFIER);
      $setuphold(posedge CP &&& EX , negedge TE, `CBUFLHSP_TE_CP_SETUP, `CBUFLHSP_TE_CP_HOLD, NOTIFIER);
      $setuphold(posedge CP &&& TEX , posedge E, `CBUFLHSP_E_CP_SETUP, `CBUFLHSP_E_CP_HOLD, NOTIFIER);
      $setuphold(posedge CP &&& TEX , negedge E, `CBUFLHSP_E_CP_SETUP, `CBUFLHSP_E_CP_HOLD, NOTIFIER);
      $width(negedge CP, `CBUFLHSP_CP_PWL, 0, NOTIFIER);


	endspecify

`endif

endmodule // CBUFLHSP

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
 
//  START
// CELL CBUFLHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define CBUFLHSX4_CP_F_G_F 0.1
`define CBUFLHSX4_CP_R_G_R 0.1
`define CBUFLHSX4_E_CP_HOLD 0.1
`define CBUFLHSX4_E_CP_SETUP 0.1
`define CBUFLHSX4_TE_CP_HOLD 0.1
`define CBUFLHSX4_TE_CP_SETUP 0.1
`define CBUFLHSX4_CP_PWL 0.1


module CBUFLHSX4 (G, CP, E, TE );

	output G;
	input CP;
	input E;
	input TE;

   reg NOTIFIER;

	or    u0 (INTERNAL1, E, TE) ;
	U_LD_N_NOTI u1 (IQ, INTERNAL1, CP , NOTIFIER) ;
	and    u2 (INTERNAL2, IQ, CP) ;
	buf    u3 (G, INTERNAL2) ;


`ifdef functional
`else
   not  (TEX, TE);
   not  (EX, E);

	specify

		(CP +=> G) = (`CBUFLHSX4_CP_R_G_R,`CBUFLHSX4_CP_F_G_F);
      $setuphold(posedge CP &&& EX , posedge TE, `CBUFLHSX4_TE_CP_SETUP, `CBUFLHSX4_TE_CP_HOLD, NOTIFIER);
      $setuphold(posedge CP &&& EX , negedge TE, `CBUFLHSX4_TE_CP_SETUP, `CBUFLHSX4_TE_CP_HOLD, NOTIFIER);
      $setuphold(posedge CP &&& TEX , posedge E, `CBUFLHSX4_E_CP_SETUP, `CBUFLHSX4_E_CP_HOLD, NOTIFIER);
      $setuphold(posedge CP &&& TEX , negedge E, `CBUFLHSX4_E_CP_SETUP, `CBUFLHSX4_E_CP_HOLD, NOTIFIER);
      $width(negedge CP, `CBUFLHSX4_CP_PWL, 0, NOTIFIER);


	endspecify

`endif

endmodule // CBUFLHSX4

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
 
//  START
// CELL DC24HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define DC24HS_A1_F_Z3N_R 0.1
`define DC24HS_A1_R_Z3N_F 0.1
`define DC24HS_A0_F_Z3N_R 0.1
`define DC24HS_A0_R_Z3N_F 0.1
`define DC24HS_A1_F_Z2N_R 0.1
`define DC24HS_A1_R_Z2N_F 0.1
`define DC24HS_A0_F_Z2N_F 0.1
`define DC24HS_A0_R_Z2N_R 0.1
`define DC24HS_A1_F_Z1N_F 0.1
`define DC24HS_A1_R_Z1N_R 0.1
`define DC24HS_A0_F_Z1N_R 0.1
`define DC24HS_A0_R_Z1N_F 0.1
`define DC24HS_A1_F_Z0N_F 0.1
`define DC24HS_A1_R_Z0N_R 0.1
`define DC24HS_A0_F_Z0N_F 0.1
`define DC24HS_A0_R_Z0N_R 0.1

module DC24HS (Z0N, Z1N, Z2N, Z3N, A0, A1);

   output Z0N;
   output Z1N;
   output Z2N;
   output Z3N;
   input A0;
   input A1;


   or  u0 (Z0N, A0, A1);
   nand  u1 (Z1N, A0, A1X);
   not  u2 (A1X, A1);
   nand  u3 (Z2N, A0X, A1);
   not  u4 (A0X, A0);
   nand  u5 (Z3N, A0, A1);


`ifdef functional
`else
   specify

      (A1 -=> Z3N) = (`DC24HS_A1_F_Z3N_R,`DC24HS_A1_R_Z3N_F);
      (A0 -=> Z3N) = (`DC24HS_A0_F_Z3N_R,`DC24HS_A0_R_Z3N_F);
      (A1 -=> Z2N) = (`DC24HS_A1_F_Z2N_R,`DC24HS_A1_R_Z2N_F);
      (A0 +=> Z2N) = (`DC24HS_A0_R_Z2N_R,`DC24HS_A0_F_Z2N_F);
      (A1 +=> Z1N) = (`DC24HS_A1_R_Z1N_R,`DC24HS_A1_F_Z1N_F);
      (A0 -=> Z1N) = (`DC24HS_A0_F_Z1N_R,`DC24HS_A0_R_Z1N_F);
      (A1 +=> Z0N) = (`DC24HS_A1_R_Z0N_R,`DC24HS_A1_F_Z0N_F);
      (A0 +=> Z0N) = (`DC24HS_A0_R_Z0N_R,`DC24HS_A0_F_Z0N_F);

   endspecify
`endif


endmodule // DC24HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:25 and Version :1.1 //
 
//  START 
// CELL DC38HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define DC38HS_A2_F_Z7N_R 0.1
`define DC38HS_A2_R_Z7N_F 0.1
`define DC38HS_A1_F_Z7N_R 0.1
`define DC38HS_A1_R_Z7N_F 0.1
`define DC38HS_A0_F_Z7N_R 0.1
`define DC38HS_A0_R_Z7N_F 0.1
`define DC38HS_A2_F_Z6N_R 0.1
`define DC38HS_A2_R_Z6N_F 0.1
`define DC38HS_A1_F_Z6N_R 0.1
`define DC38HS_A1_R_Z6N_F 0.1
`define DC38HS_A0_F_Z6N_F 0.1
`define DC38HS_A0_R_Z6N_R 0.1
`define DC38HS_A2_F_Z5N_R 0.1
`define DC38HS_A2_R_Z5N_F 0.1
`define DC38HS_A1_F_Z5N_F 0.1
`define DC38HS_A1_R_Z5N_R 0.1
`define DC38HS_A0_F_Z5N_R 0.1
`define DC38HS_A0_R_Z5N_F 0.1
`define DC38HS_A2_F_Z4N_R 0.1
`define DC38HS_A2_R_Z4N_F 0.1
`define DC38HS_A1_F_Z4N_F 0.1
`define DC38HS_A1_R_Z4N_R 0.1
`define DC38HS_A0_F_Z4N_F 0.1
`define DC38HS_A0_R_Z4N_R 0.1
`define DC38HS_A2_F_Z3N_F 0.1
`define DC38HS_A2_R_Z3N_R 0.1
`define DC38HS_A1_F_Z3N_R 0.1
`define DC38HS_A1_R_Z3N_F 0.1
`define DC38HS_A0_F_Z3N_R 0.1
`define DC38HS_A0_R_Z3N_F 0.1
`define DC38HS_A2_F_Z2N_F 0.1
`define DC38HS_A2_R_Z2N_R 0.1
`define DC38HS_A1_F_Z2N_R 0.1
`define DC38HS_A1_R_Z2N_F 0.1
`define DC38HS_A0_F_Z2N_F 0.1
`define DC38HS_A0_R_Z2N_R 0.1
`define DC38HS_A2_F_Z1N_F 0.1
`define DC38HS_A2_R_Z1N_R 0.1
`define DC38HS_A1_F_Z1N_F 0.1
`define DC38HS_A1_R_Z1N_R 0.1
`define DC38HS_A0_F_Z1N_R 0.1
`define DC38HS_A0_R_Z1N_F 0.1
`define DC38HS_A2_F_Z0N_F 0.1
`define DC38HS_A2_R_Z0N_R 0.1
`define DC38HS_A1_F_Z0N_F 0.1
`define DC38HS_A1_R_Z0N_R 0.1
`define DC38HS_A0_F_Z0N_F 0.1
`define DC38HS_A0_R_Z0N_R 0.1

module DC38HS (Z0N, Z1N, Z2N, Z3N, Z4N, Z5N, Z6N, Z7N, A0, A1, A2);

   output Z0N;
   output Z1N;
   output Z2N;
   output Z3N;
   output Z4N;
   output Z5N;
   output Z6N;
   output Z7N;
   input A0;
   input A1;
   input A2;


   or  u0 (Z0N, A0, A1, A2);
   or  u1 (Z1N, A0X, A1, A2);
   not  u2 (A0X, A0);
   or  u3 (Z2N, A0, A1X, A2);
   not  u4 (A1X, A1);
   nand  u5 (Z3N, A0, A1, A2X);
   not  u6 (A2X, A2);
   or  u7 (Z4N, A0, A1, A2X);
   nand  u8 (Z5N, A0, A1X, A2);
   nand  u9 (Z6N, A0X, A1, A2);
   nand  u10 (Z7N, A0, A1, A2);


`ifdef functional
`else
   specify

      (A2 -=> Z7N) = (`DC38HS_A2_F_Z7N_R,`DC38HS_A2_R_Z7N_F);
      (A1 -=> Z7N) = (`DC38HS_A1_F_Z7N_R,`DC38HS_A1_R_Z7N_F);
      (A0 -=> Z7N) = (`DC38HS_A0_F_Z7N_R,`DC38HS_A0_R_Z7N_F);
      (A2 -=> Z6N) = (`DC38HS_A2_F_Z6N_R,`DC38HS_A2_R_Z6N_F);
      (A1 -=> Z6N) = (`DC38HS_A1_F_Z6N_R,`DC38HS_A1_R_Z6N_F);
      (A0 +=> Z6N) = (`DC38HS_A0_R_Z6N_R,`DC38HS_A0_F_Z6N_F);
      (A2 -=> Z5N) = (`DC38HS_A2_F_Z5N_R,`DC38HS_A2_R_Z5N_F);
      (A1 +=> Z5N) = (`DC38HS_A1_R_Z5N_R,`DC38HS_A1_F_Z5N_F);
      (A0 -=> Z5N) = (`DC38HS_A0_F_Z5N_R,`DC38HS_A0_R_Z5N_F);
      (A2 -=> Z4N) = (`DC38HS_A2_F_Z4N_R,`DC38HS_A2_R_Z4N_F);
      (A1 +=> Z4N) = (`DC38HS_A1_R_Z4N_R,`DC38HS_A1_F_Z4N_F);
      (A0 +=> Z4N) = (`DC38HS_A0_R_Z4N_R,`DC38HS_A0_F_Z4N_F);
      (A2 +=> Z3N) = (`DC38HS_A2_R_Z3N_R,`DC38HS_A2_F_Z3N_F);
      (A1 -=> Z3N) = (`DC38HS_A1_F_Z3N_R,`DC38HS_A1_R_Z3N_F);
      (A0 -=> Z3N) = (`DC38HS_A0_F_Z3N_R,`DC38HS_A0_R_Z3N_F);
      (A2 +=> Z2N) = (`DC38HS_A2_R_Z2N_R,`DC38HS_A2_F_Z2N_F);
      (A1 -=> Z2N) = (`DC38HS_A1_F_Z2N_R,`DC38HS_A1_R_Z2N_F);
      (A0 +=> Z2N) = (`DC38HS_A0_R_Z2N_R,`DC38HS_A0_F_Z2N_F);
      (A2 +=> Z1N) = (`DC38HS_A2_R_Z1N_R,`DC38HS_A2_F_Z1N_F);
      (A1 +=> Z1N) = (`DC38HS_A1_R_Z1N_R,`DC38HS_A1_F_Z1N_F);
      (A0 -=> Z1N) = (`DC38HS_A0_F_Z1N_R,`DC38HS_A0_R_Z1N_F);
      (A2 +=> Z0N) = (`DC38HS_A2_R_Z0N_R,`DC38HS_A2_F_Z0N_F);
      (A1 +=> Z0N) = (`DC38HS_A1_R_Z0N_R,`DC38HS_A1_F_Z0N_F);
      (A0 +=> Z0N) = (`DC38HS_A0_R_Z0N_R,`DC38HS_A0_F_Z0N_F);

   endspecify
`endif


endmodule // DC38HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:29 and Version :1.1 //
 
//  START 
// CELL DE24HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define DE24HS_A1_F_Z3N_R 0.1
`define DE24HS_A1_R_Z3N_F 0.1
`define DE24HS_A0_F_Z3N_R 0.1
`define DE24HS_A0_R_Z3N_F 0.1
`define DE24HS_EN_F_Z3N_F 0.1
`define DE24HS_EN_R_Z3N_R 0.1
`define DE24HS_A1_F_Z2N_R 0.1
`define DE24HS_A1_R_Z2N_F 0.1
`define DE24HS_A0_F_Z2N_F 0.1
`define DE24HS_A0_R_Z2N_R 0.1
`define DE24HS_EN_F_Z2N_F 0.1
`define DE24HS_EN_R_Z2N_R 0.1
`define DE24HS_A1_F_Z1N_F 0.1
`define DE24HS_A1_R_Z1N_R 0.1
`define DE24HS_A0_F_Z1N_R 0.1
`define DE24HS_A0_R_Z1N_F 0.1
`define DE24HS_EN_F_Z1N_F 0.1
`define DE24HS_EN_R_Z1N_R 0.1
`define DE24HS_A1_F_Z0N_F 0.1
`define DE24HS_A1_R_Z0N_R 0.1
`define DE24HS_A0_F_Z0N_F 0.1
`define DE24HS_A0_R_Z0N_R 0.1
`define DE24HS_EN_F_Z0N_F 0.1
`define DE24HS_EN_R_Z0N_R 0.1

module DE24HS (Z0N, Z1N, Z2N, Z3N, A0, A1, EN);

   output Z0N;
   output Z1N;
   output Z2N;
   output Z3N;
   input EN;
   input A0;
   input A1;


   or  u0 (Z0N, A0, A1, EN);
   or  u1 (Z1N, A0X, A1, EN);
   not  u2 (A0X, A0);
   or  u3 (Z2N, A0, A1X, EN);
   not  u4 (A1X, A1);
   nand  u5 (Z3N, A0, A1, ENX);
   not  u6 (ENX, EN);


`ifdef functional
`else
   specify

      (A1 -=> Z3N) = (`DE24HS_A1_F_Z3N_R,`DE24HS_A1_R_Z3N_F);
      (A0 -=> Z3N) = (`DE24HS_A0_F_Z3N_R,`DE24HS_A0_R_Z3N_F);
      (EN +=> Z3N) = (`DE24HS_EN_R_Z3N_R,`DE24HS_EN_F_Z3N_F);
      (A1 -=> Z2N) = (`DE24HS_A1_F_Z2N_R,`DE24HS_A1_R_Z2N_F);
      (A0 +=> Z2N) = (`DE24HS_A0_R_Z2N_R,`DE24HS_A0_F_Z2N_F);
      (EN +=> Z2N) = (`DE24HS_EN_R_Z2N_R,`DE24HS_EN_F_Z2N_F);
      (A1 +=> Z1N) = (`DE24HS_A1_R_Z1N_R,`DE24HS_A1_F_Z1N_F);
      (A0 -=> Z1N) = (`DE24HS_A0_F_Z1N_R,`DE24HS_A0_R_Z1N_F);
      (EN +=> Z1N) = (`DE24HS_EN_R_Z1N_R,`DE24HS_EN_F_Z1N_F);
      (A1 +=> Z0N) = (`DE24HS_A1_R_Z0N_R,`DE24HS_A1_F_Z0N_F);
      (A0 +=> Z0N) = (`DE24HS_A0_R_Z0N_R,`DE24HS_A0_F_Z0N_F);
      (EN +=> Z0N) = (`DE24HS_EN_R_Z0N_R,`DE24HS_EN_F_Z0N_F);

   endspecify
`endif


endmodule // DE24HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:32 and Version :1.1 //
 
//  START 
// CELL ENHSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ENHSX05_B_F_Z_F 0.1
`define ENHSX05_B_R_Z_R 0.1
`define ENHSX05_B_F_Z_R 0.1
`define ENHSX05_B_R_Z_F 0.1
`define ENHSX05_A_F_Z_F 0.1
`define ENHSX05_A_R_Z_R 0.1
`define ENHSX05_A_F_Z_R 0.1
`define ENHSX05_A_R_Z_F 0.1

module ENHSX05 (Z, A, B);

   output Z;
   input A;
   input B;


   xnor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      if (A) (B +=> Z) = (`ENHSX05_B_R_Z_R,`ENHSX05_B_F_Z_F);
      if (!A) (B -=> Z) = (`ENHSX05_B_F_Z_R,`ENHSX05_B_R_Z_F);
      if (B) (A +=> Z) = (`ENHSX05_A_R_Z_R,`ENHSX05_A_F_Z_F);
      if (!B) (A -=> Z) = (`ENHSX05_A_F_Z_R,`ENHSX05_A_R_Z_F);

   endspecify
`endif


endmodule // ENHSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:41 and Version :1.1 //
 
//  START 
// CELL ENHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ENHS_B_F_Z_F 0.1
`define ENHS_B_R_Z_R 0.1
`define ENHS_B_F_Z_R 0.1
`define ENHS_B_R_Z_F 0.1
`define ENHS_A_F_Z_F 0.1
`define ENHS_A_R_Z_R 0.1
`define ENHS_A_F_Z_R 0.1
`define ENHS_A_R_Z_F 0.1

module ENHS (Z, A, B);

   output Z;
   input A;
   input B;


   xnor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      if (A) (B +=> Z) = (`ENHS_B_R_Z_R,`ENHS_B_F_Z_F);
      if (!A) (B -=> Z) = (`ENHS_B_F_Z_R,`ENHS_B_R_Z_F);
      if (B) (A +=> Z) = (`ENHS_A_R_Z_R,`ENHS_A_F_Z_F);
      if (!B) (A -=> Z) = (`ENHS_A_F_Z_R,`ENHS_A_R_Z_F);

   endspecify
`endif


endmodule // ENHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:41 and Version :1.1 //
 
//  START 
// CELL ENHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ENHSP_B_F_Z_F 0.1
`define ENHSP_B_R_Z_R 0.1
`define ENHSP_B_F_Z_R 0.1
`define ENHSP_B_R_Z_F 0.1
`define ENHSP_A_F_Z_F 0.1
`define ENHSP_A_R_Z_R 0.1
`define ENHSP_A_F_Z_R 0.1
`define ENHSP_A_R_Z_F 0.1

module ENHSP (Z, A, B);

   output Z;
   input A;
   input B;


   xnor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      if (A) (B +=> Z) = (`ENHSP_B_R_Z_R,`ENHSP_B_F_Z_F);
      if (!A) (B -=> Z) = (`ENHSP_B_F_Z_R,`ENHSP_B_R_Z_F);
      if (B) (A +=> Z) = (`ENHSP_A_R_Z_R,`ENHSP_A_F_Z_F);
      if (!B) (A -=> Z) = (`ENHSP_A_F_Z_R,`ENHSP_A_R_Z_F);

   endspecify
`endif


endmodule // ENHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:41 and Version :1.1 //
 
//  START 
// CELL ENHSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ENHSX3_B_F_Z_F 0.1
`define ENHSX3_B_R_Z_R 0.1
`define ENHSX3_B_F_Z_R 0.1
`define ENHSX3_B_R_Z_F 0.1
`define ENHSX3_A_F_Z_F 0.1
`define ENHSX3_A_R_Z_R 0.1
`define ENHSX3_A_F_Z_R 0.1
`define ENHSX3_A_R_Z_F 0.1

module ENHSX3 (Z, A, B);

   output Z;
   input A;
   input B;


   xnor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      if (A) (B +=> Z) = (`ENHSX3_B_R_Z_R,`ENHSX3_B_F_Z_F);
      if (!A) (B -=> Z) = (`ENHSX3_B_F_Z_R,`ENHSX3_B_R_Z_F);
      if (B) (A +=> Z) = (`ENHSX3_A_R_Z_R,`ENHSX3_A_F_Z_F);
      if (!B) (A -=> Z) = (`ENHSX3_A_F_Z_R,`ENHSX3_A_R_Z_F);

   endspecify
`endif


endmodule // ENHSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:41 and Version :1.1 //
 
//  START 
// CELL ENHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ENHSX4_B_F_Z_F 0.1
`define ENHSX4_B_R_Z_R 0.1
`define ENHSX4_B_F_Z_R 0.1
`define ENHSX4_B_R_Z_F 0.1
`define ENHSX4_A_F_Z_F 0.1
`define ENHSX4_A_R_Z_R 0.1
`define ENHSX4_A_F_Z_R 0.1
`define ENHSX4_A_R_Z_F 0.1

module ENHSX4 (Z, A, B);

   output Z;
   input A;
   input B;


   xnor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      if (A) (B +=> Z) = (`ENHSX4_B_R_Z_R,`ENHSX4_B_F_Z_F);
      if (!A) (B -=> Z) = (`ENHSX4_B_F_Z_R,`ENHSX4_B_R_Z_F);
      if (B) (A +=> Z) = (`ENHSX4_A_R_Z_R,`ENHSX4_A_F_Z_F);
      if (!B) (A -=> Z) = (`ENHSX4_A_F_Z_R,`ENHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // ENHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:41 and Version :1.1 //
 
//  START 
// CELL F_ENHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_ENHSP_B_F_Z_F 0.1
`define F_ENHSP_B_R_Z_R 0.1
`define F_ENHSP_B_F_Z_R 0.1
`define F_ENHSP_B_R_Z_F 0.1
`define F_ENHSP_A_F_Z_F 0.1
`define F_ENHSP_A_R_Z_R 0.1
`define F_ENHSP_A_F_Z_R 0.1
`define F_ENHSP_A_R_Z_F 0.1

module F_ENHSP (Z, A, B);

   output Z;
   input A;
   input B;


   xnor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      if (A) (B +=> Z) = (`F_ENHSP_B_R_Z_R,`F_ENHSP_B_F_Z_F);
      if (!A) (B -=> Z) = (`F_ENHSP_B_F_Z_R,`F_ENHSP_B_R_Z_F);
      if (B) (A +=> Z) = (`F_ENHSP_A_R_Z_R,`F_ENHSP_A_F_Z_F);
      if (!B) (A -=> Z) = (`F_ENHSP_A_F_Z_R,`F_ENHSP_A_R_Z_F);

   endspecify
`endif


endmodule // F_ENHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:41 and Version :1.1 //
 
//  START 
// CELL F_ENHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_ENHSX4_B_F_Z_F 0.1
`define F_ENHSX4_B_R_Z_R 0.1
`define F_ENHSX4_B_F_Z_R 0.1
`define F_ENHSX4_B_R_Z_F 0.1
`define F_ENHSX4_A_F_Z_F 0.1
`define F_ENHSX4_A_R_Z_R 0.1
`define F_ENHSX4_A_F_Z_R 0.1
`define F_ENHSX4_A_R_Z_F 0.1

module F_ENHSX4 (Z, A, B);

   output Z;
   input A;
   input B;


   xnor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      if (A) (B +=> Z) = (`F_ENHSX4_B_R_Z_R,`F_ENHSX4_B_F_Z_F);
      if (!A) (B -=> Z) = (`F_ENHSX4_B_F_Z_R,`F_ENHSX4_B_R_Z_F);
      if (B) (A +=> Z) = (`F_ENHSX4_A_R_Z_R,`F_ENHSX4_A_F_Z_F);
      if (!B) (A -=> Z) = (`F_ENHSX4_A_F_Z_R,`F_ENHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // F_ENHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:41 and Version :1.1 //
 
//  START 
// CELL EN3HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define EN3HSX05_C_F_Z_R 0.1
`define EN3HSX05_C_R_Z_F 0.1
`define EN3HSX05_C_F_Z_F 0.1
`define EN3HSX05_C_R_Z_R 0.1
`define EN3HSX05_B_F_Z_R 0.1
`define EN3HSX05_B_R_Z_F 0.1
`define EN3HSX05_B_F_Z_F 0.1
`define EN3HSX05_B_R_Z_R 0.1
`define EN3HSX05_A_F_Z_R 0.1
`define EN3HSX05_A_R_Z_F 0.1
`define EN3HSX05_A_F_Z_F 0.1
`define EN3HSX05_A_R_Z_R 0.1

module EN3HSX05 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   xnor  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      if (A && B || !A && !B) (C -=> Z) = (`EN3HSX05_C_F_Z_R,`EN3HSX05_C_R_Z_F);
      if (!A && B || A && !B) (C +=> Z) = (`EN3HSX05_C_R_Z_R,`EN3HSX05_C_F_Z_F);
      if (A && C || !A && !C) (B -=> Z) = (`EN3HSX05_B_F_Z_R,`EN3HSX05_B_R_Z_F);
      if (!A && C || A && !C) (B +=> Z) = (`EN3HSX05_B_R_Z_R,`EN3HSX05_B_F_Z_F);
      if (B && C || !B && !C) (A -=> Z) = (`EN3HSX05_A_F_Z_R,`EN3HSX05_A_R_Z_F);
      if (!B && C || B && !C) (A +=> Z) = (`EN3HSX05_A_R_Z_R,`EN3HSX05_A_F_Z_F);

   endspecify
`endif


endmodule // EN3HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:41 and Version :1.1 //
 
//  START 
// CELL EN3HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define EN3HS_C_F_Z_R 0.1
`define EN3HS_C_R_Z_F 0.1
`define EN3HS_C_F_Z_F 0.1
`define EN3HS_C_R_Z_R 0.1
`define EN3HS_B_F_Z_R 0.1
`define EN3HS_B_R_Z_F 0.1
`define EN3HS_B_F_Z_F 0.1
`define EN3HS_B_R_Z_R 0.1
`define EN3HS_A_F_Z_R 0.1
`define EN3HS_A_R_Z_F 0.1
`define EN3HS_A_F_Z_F 0.1
`define EN3HS_A_R_Z_R 0.1

module EN3HS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   xnor  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      if (A && B || !A && !B) (C -=> Z) = (`EN3HS_C_F_Z_R,`EN3HS_C_R_Z_F);
      if (!A && B || A && !B) (C +=> Z) = (`EN3HS_C_R_Z_R,`EN3HS_C_F_Z_F);
      if (A && C || !A && !C) (B -=> Z) = (`EN3HS_B_F_Z_R,`EN3HS_B_R_Z_F);
      if (!A && C || A && !C) (B +=> Z) = (`EN3HS_B_R_Z_R,`EN3HS_B_F_Z_F);
      if (B && C || !B && !C) (A -=> Z) = (`EN3HS_A_F_Z_R,`EN3HS_A_R_Z_F);
      if (!B && C || B && !C) (A +=> Z) = (`EN3HS_A_R_Z_R,`EN3HS_A_F_Z_F);

   endspecify
`endif


endmodule // EN3HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:41 and Version :1.1 //
 
//  START 
// CELL EN3HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define EN3HSP_C_F_Z_R 0.1
`define EN3HSP_C_R_Z_F 0.1
`define EN3HSP_C_F_Z_F 0.1
`define EN3HSP_C_R_Z_R 0.1
`define EN3HSP_B_F_Z_R 0.1
`define EN3HSP_B_R_Z_F 0.1
`define EN3HSP_B_F_Z_F 0.1
`define EN3HSP_B_R_Z_R 0.1
`define EN3HSP_A_F_Z_R 0.1
`define EN3HSP_A_R_Z_F 0.1
`define EN3HSP_A_F_Z_F 0.1
`define EN3HSP_A_R_Z_R 0.1

module EN3HSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   xnor  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      if (A && B || !A && !B) (C -=> Z) = (`EN3HSP_C_F_Z_R,`EN3HSP_C_R_Z_F);
      if (!A && B || A && !B) (C +=> Z) = (`EN3HSP_C_R_Z_R,`EN3HSP_C_F_Z_F);
      if (A && C || !A && !C) (B -=> Z) = (`EN3HSP_B_F_Z_R,`EN3HSP_B_R_Z_F);
      if (!A && C || A && !C) (B +=> Z) = (`EN3HSP_B_R_Z_R,`EN3HSP_B_F_Z_F);
      if (B && C || !B && !C) (A -=> Z) = (`EN3HSP_A_F_Z_R,`EN3HSP_A_R_Z_F);
      if (!B && C || B && !C) (A +=> Z) = (`EN3HSP_A_R_Z_R,`EN3HSP_A_F_Z_F);

   endspecify
`endif


endmodule // EN3HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:41 and Version :1.1 //
 
//  START 
// CELL EN3HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define EN3HSX4_C_F_Z_R 0.1
`define EN3HSX4_C_R_Z_F 0.1
`define EN3HSX4_C_F_Z_F 0.1
`define EN3HSX4_C_R_Z_R 0.1
`define EN3HSX4_B_F_Z_R 0.1
`define EN3HSX4_B_R_Z_F 0.1
`define EN3HSX4_B_F_Z_F 0.1
`define EN3HSX4_B_R_Z_R 0.1
`define EN3HSX4_A_F_Z_R 0.1
`define EN3HSX4_A_R_Z_F 0.1
`define EN3HSX4_A_F_Z_F 0.1
`define EN3HSX4_A_R_Z_R 0.1

module EN3HSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   xnor  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      if (A && B || !A && !B) (C -=> Z) = (`EN3HSX4_C_F_Z_R,`EN3HSX4_C_R_Z_F);
      if (!A && B || A && !B) (C +=> Z) = (`EN3HSX4_C_R_Z_R,`EN3HSX4_C_F_Z_F);
      if (A && C || !A && !C) (B -=> Z) = (`EN3HSX4_B_F_Z_R,`EN3HSX4_B_R_Z_F);
      if (!A && C || A && !C) (B +=> Z) = (`EN3HSX4_B_R_Z_R,`EN3HSX4_B_F_Z_F);
      if (B && C || !B && !C) (A -=> Z) = (`EN3HSX4_A_F_Z_R,`EN3HSX4_A_R_Z_F);
      if (!B && C || B && !C) (A +=> Z) = (`EN3HSX4_A_R_Z_R,`EN3HSX4_A_F_Z_F);

   endspecify
`endif


endmodule // EN3HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:41 and Version :1.1 //
 
//  START 
// CELL F_EN3HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_EN3HSP_C_F_Z_R 0.1
`define F_EN3HSP_C_R_Z_F 0.1
`define F_EN3HSP_C_F_Z_F 0.1
`define F_EN3HSP_C_R_Z_R 0.1
`define F_EN3HSP_B_F_Z_R 0.1
`define F_EN3HSP_B_R_Z_F 0.1
`define F_EN3HSP_B_F_Z_F 0.1
`define F_EN3HSP_B_R_Z_R 0.1
`define F_EN3HSP_A_F_Z_R 0.1
`define F_EN3HSP_A_R_Z_F 0.1
`define F_EN3HSP_A_F_Z_F 0.1
`define F_EN3HSP_A_R_Z_R 0.1

module F_EN3HSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   xnor  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      if (A && B || !A && !B) (C -=> Z) = (`F_EN3HSP_C_F_Z_R,`F_EN3HSP_C_R_Z_F);
      if (!A && B || A && !B) (C +=> Z) = (`F_EN3HSP_C_R_Z_R,`F_EN3HSP_C_F_Z_F);
      if (A && C || !A && !C) (B -=> Z) = (`F_EN3HSP_B_F_Z_R,`F_EN3HSP_B_R_Z_F);
      if (!A && C || A && !C) (B +=> Z) = (`F_EN3HSP_B_R_Z_R,`F_EN3HSP_B_F_Z_F);
      if (B && C || !B && !C) (A -=> Z) = (`F_EN3HSP_A_F_Z_R,`F_EN3HSP_A_R_Z_F);
      if (!B && C || B && !C) (A +=> Z) = (`F_EN3HSP_A_R_Z_R,`F_EN3HSP_A_F_Z_F);

   endspecify
`endif


endmodule // F_EN3HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:41 and Version :1.1 //
 
//  START 
// CELL F_EN3HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_EN3HSX4_C_F_Z_R 0.1
`define F_EN3HSX4_C_R_Z_F 0.1
`define F_EN3HSX4_C_F_Z_F 0.1
`define F_EN3HSX4_C_R_Z_R 0.1
`define F_EN3HSX4_B_F_Z_R 0.1
`define F_EN3HSX4_B_R_Z_F 0.1
`define F_EN3HSX4_B_F_Z_F 0.1
`define F_EN3HSX4_B_R_Z_R 0.1
`define F_EN3HSX4_A_F_Z_R 0.1
`define F_EN3HSX4_A_R_Z_F 0.1
`define F_EN3HSX4_A_F_Z_F 0.1
`define F_EN3HSX4_A_R_Z_R 0.1

module F_EN3HSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   xnor  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      if (A && B || !A && !B) (C -=> Z) = (`F_EN3HSX4_C_F_Z_R,`F_EN3HSX4_C_R_Z_F);
      if (!A && B || A && !B) (C +=> Z) = (`F_EN3HSX4_C_R_Z_R,`F_EN3HSX4_C_F_Z_F);
      if (A && C || !A && !C) (B -=> Z) = (`F_EN3HSX4_B_F_Z_R,`F_EN3HSX4_B_R_Z_F);
      if (!A && C || A && !C) (B +=> Z) = (`F_EN3HSX4_B_R_Z_R,`F_EN3HSX4_B_F_Z_F);
      if (B && C || !B && !C) (A -=> Z) = (`F_EN3HSX4_A_F_Z_R,`F_EN3HSX4_A_R_Z_F);
      if (!B && C || B && !C) (A +=> Z) = (`F_EN3HSX4_A_R_Z_R,`F_EN3HSX4_A_F_Z_F);

   endspecify
`endif


endmodule // F_EN3HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:41 and Version :1.1 //
 
//  START 
// CELL EOHSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define EOHSX05_B_F_Z_R 0.1
`define EOHSX05_B_R_Z_F 0.1
`define EOHSX05_B_F_Z_F 0.1
`define EOHSX05_B_R_Z_R 0.1
`define EOHSX05_A_F_Z_R 0.1
`define EOHSX05_A_R_Z_F 0.1
`define EOHSX05_A_F_Z_F 0.1
`define EOHSX05_A_R_Z_R 0.1

module EOHSX05 (Z, A, B);

   output Z;
   input A;
   input B;


   xor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      if (A) (B -=> Z) = (`EOHSX05_B_F_Z_R,`EOHSX05_B_R_Z_F);
      if (!A) (B +=> Z) = (`EOHSX05_B_R_Z_R,`EOHSX05_B_F_Z_F);
      if (B) (A -=> Z) = (`EOHSX05_A_F_Z_R,`EOHSX05_A_R_Z_F);
      if (!B) (A +=> Z) = (`EOHSX05_A_R_Z_R,`EOHSX05_A_F_Z_F);

   endspecify
`endif


endmodule // EOHSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:47 and Version :1.1 //
 
//  START 
// CELL EOHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define EOHS_B_F_Z_R 0.1
`define EOHS_B_R_Z_F 0.1
`define EOHS_B_F_Z_F 0.1
`define EOHS_B_R_Z_R 0.1
`define EOHS_A_F_Z_R 0.1
`define EOHS_A_R_Z_F 0.1
`define EOHS_A_F_Z_F 0.1
`define EOHS_A_R_Z_R 0.1

module EOHS (Z, A, B);

   output Z;
   input A;
   input B;


   xor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      if (A) (B -=> Z) = (`EOHS_B_F_Z_R,`EOHS_B_R_Z_F);
      if (!A) (B +=> Z) = (`EOHS_B_R_Z_R,`EOHS_B_F_Z_F);
      if (B) (A -=> Z) = (`EOHS_A_F_Z_R,`EOHS_A_R_Z_F);
      if (!B) (A +=> Z) = (`EOHS_A_R_Z_R,`EOHS_A_F_Z_F);

   endspecify
`endif


endmodule // EOHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:47 and Version :1.1 //
 
//  START 
// CELL EOHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define EOHSP_B_F_Z_R 0.1
`define EOHSP_B_R_Z_F 0.1
`define EOHSP_B_F_Z_F 0.1
`define EOHSP_B_R_Z_R 0.1
`define EOHSP_A_F_Z_R 0.1
`define EOHSP_A_R_Z_F 0.1
`define EOHSP_A_F_Z_F 0.1
`define EOHSP_A_R_Z_R 0.1

module EOHSP (Z, A, B);

   output Z;
   input A;
   input B;


   xor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      if (A) (B -=> Z) = (`EOHSP_B_F_Z_R,`EOHSP_B_R_Z_F);
      if (!A) (B +=> Z) = (`EOHSP_B_R_Z_R,`EOHSP_B_F_Z_F);
      if (B) (A -=> Z) = (`EOHSP_A_F_Z_R,`EOHSP_A_R_Z_F);
      if (!B) (A +=> Z) = (`EOHSP_A_R_Z_R,`EOHSP_A_F_Z_F);

   endspecify
`endif


endmodule // EOHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:47 and Version :1.1 //
 
//  START 
// CELL EOHSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define EOHSX3_B_F_Z_R 0.1
`define EOHSX3_B_R_Z_F 0.1
`define EOHSX3_B_F_Z_F 0.1
`define EOHSX3_B_R_Z_R 0.1
`define EOHSX3_A_F_Z_R 0.1
`define EOHSX3_A_R_Z_F 0.1
`define EOHSX3_A_F_Z_F 0.1
`define EOHSX3_A_R_Z_R 0.1

module EOHSX3 (Z, A, B);

   output Z;
   input A;
   input B;


   xor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      if (A) (B -=> Z) = (`EOHSX3_B_F_Z_R,`EOHSX3_B_R_Z_F);
      if (!A) (B +=> Z) = (`EOHSX3_B_R_Z_R,`EOHSX3_B_F_Z_F);
      if (B) (A -=> Z) = (`EOHSX3_A_F_Z_R,`EOHSX3_A_R_Z_F);
      if (!B) (A +=> Z) = (`EOHSX3_A_R_Z_R,`EOHSX3_A_F_Z_F);

   endspecify
`endif


endmodule // EOHSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:47 and Version :1.1 //
 
//  START 
// CELL EOHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define EOHSX4_B_F_Z_R 0.1
`define EOHSX4_B_R_Z_F 0.1
`define EOHSX4_B_F_Z_F 0.1
`define EOHSX4_B_R_Z_R 0.1
`define EOHSX4_A_F_Z_R 0.1
`define EOHSX4_A_R_Z_F 0.1
`define EOHSX4_A_F_Z_F 0.1
`define EOHSX4_A_R_Z_R 0.1

module EOHSX4 (Z, A, B);

   output Z;
   input A;
   input B;


   xor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      if (A) (B -=> Z) = (`EOHSX4_B_F_Z_R,`EOHSX4_B_R_Z_F);
      if (!A) (B +=> Z) = (`EOHSX4_B_R_Z_R,`EOHSX4_B_F_Z_F);
      if (B) (A -=> Z) = (`EOHSX4_A_F_Z_R,`EOHSX4_A_R_Z_F);
      if (!B) (A +=> Z) = (`EOHSX4_A_R_Z_R,`EOHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // EOHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:47 and Version :1.1 //
 
//  START 
// CELL F_EOHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_EOHS_B_F_Z_R 0.1
`define F_EOHS_B_R_Z_F 0.1
`define F_EOHS_B_F_Z_F 0.1
`define F_EOHS_B_R_Z_R 0.1
`define F_EOHS_A_F_Z_R 0.1
`define F_EOHS_A_R_Z_F 0.1
`define F_EOHS_A_F_Z_F 0.1
`define F_EOHS_A_R_Z_R 0.1

module F_EOHS (Z, A, B);

   output Z;
   input A;
   input B;


   xor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      if (A) (B -=> Z) = (`F_EOHS_B_F_Z_R,`F_EOHS_B_R_Z_F);
      if (!A) (B +=> Z) = (`F_EOHS_B_R_Z_R,`F_EOHS_B_F_Z_F);
      if (B) (A -=> Z) = (`F_EOHS_A_F_Z_R,`F_EOHS_A_R_Z_F);
      if (!B) (A +=> Z) = (`F_EOHS_A_R_Z_R,`F_EOHS_A_F_Z_F);

   endspecify
`endif


endmodule // F_EOHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:47 and Version :1.1 //
 
//  START 
// CELL F_EOHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_EOHSP_B_F_Z_R 0.1
`define F_EOHSP_B_R_Z_F 0.1
`define F_EOHSP_B_F_Z_F 0.1
`define F_EOHSP_B_R_Z_R 0.1
`define F_EOHSP_A_F_Z_R 0.1
`define F_EOHSP_A_R_Z_F 0.1
`define F_EOHSP_A_F_Z_F 0.1
`define F_EOHSP_A_R_Z_R 0.1

module F_EOHSP (Z, A, B);

   output Z;
   input A;
   input B;


   xor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      if (A) (B -=> Z) = (`F_EOHSP_B_F_Z_R,`F_EOHSP_B_R_Z_F);
      if (!A) (B +=> Z) = (`F_EOHSP_B_R_Z_R,`F_EOHSP_B_F_Z_F);
      if (B) (A -=> Z) = (`F_EOHSP_A_F_Z_R,`F_EOHSP_A_R_Z_F);
      if (!B) (A +=> Z) = (`F_EOHSP_A_R_Z_R,`F_EOHSP_A_F_Z_F);

   endspecify
`endif


endmodule // F_EOHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:47 and Version :1.1 //
 
//  START 
// CELL F_EOHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_EOHSX4_B_F_Z_R 0.1
`define F_EOHSX4_B_R_Z_F 0.1
`define F_EOHSX4_B_F_Z_F 0.1
`define F_EOHSX4_B_R_Z_R 0.1
`define F_EOHSX4_A_F_Z_R 0.1
`define F_EOHSX4_A_R_Z_F 0.1
`define F_EOHSX4_A_F_Z_F 0.1
`define F_EOHSX4_A_R_Z_R 0.1

module F_EOHSX4 (Z, A, B);

   output Z;
   input A;
   input B;


   xor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      if (A) (B -=> Z) = (`F_EOHSX4_B_F_Z_R,`F_EOHSX4_B_R_Z_F);
      if (!A) (B +=> Z) = (`F_EOHSX4_B_R_Z_R,`F_EOHSX4_B_F_Z_F);
      if (B) (A -=> Z) = (`F_EOHSX4_A_F_Z_R,`F_EOHSX4_A_R_Z_F);
      if (!B) (A +=> Z) = (`F_EOHSX4_A_R_Z_R,`F_EOHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // F_EOHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:47 and Version :1.1 //
 
//  START 
// CELL EO3HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define EO3HSX05_C_F_Z_F 0.1
`define EO3HSX05_C_R_Z_R 0.1
`define EO3HSX05_C_F_Z_R 0.1
`define EO3HSX05_C_R_Z_F 0.1
`define EO3HSX05_B_F_Z_F 0.1
`define EO3HSX05_B_R_Z_R 0.1
`define EO3HSX05_B_F_Z_R 0.1
`define EO3HSX05_B_R_Z_F 0.1
`define EO3HSX05_A_F_Z_F 0.1
`define EO3HSX05_A_R_Z_R 0.1
`define EO3HSX05_A_F_Z_R 0.1
`define EO3HSX05_A_R_Z_F 0.1

module EO3HSX05 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   xor  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      if (A && B || !A && !B) (C +=> Z) = (`EO3HSX05_C_R_Z_R,`EO3HSX05_C_F_Z_F);
      if (!A && B || A && !B) (C -=> Z) = (`EO3HSX05_C_F_Z_R,`EO3HSX05_C_R_Z_F);
      if (A && C || !A && !C) (B +=> Z) = (`EO3HSX05_B_R_Z_R,`EO3HSX05_B_F_Z_F);
      if (!A && C || A && !C) (B -=> Z) = (`EO3HSX05_B_F_Z_R,`EO3HSX05_B_R_Z_F);
      if (B && C || !B && !C) (A +=> Z) = (`EO3HSX05_A_R_Z_R,`EO3HSX05_A_F_Z_F);
      if (!B && C || B && !C) (A -=> Z) = (`EO3HSX05_A_F_Z_R,`EO3HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // EO3HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:47 and Version :1.1 //
 
//  START 
// CELL EO3HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define EO3HS_C_F_Z_F 0.1
`define EO3HS_C_R_Z_R 0.1
`define EO3HS_C_F_Z_R 0.1
`define EO3HS_C_R_Z_F 0.1
`define EO3HS_B_F_Z_F 0.1
`define EO3HS_B_R_Z_R 0.1
`define EO3HS_B_F_Z_R 0.1
`define EO3HS_B_R_Z_F 0.1
`define EO3HS_A_F_Z_F 0.1
`define EO3HS_A_R_Z_R 0.1
`define EO3HS_A_F_Z_R 0.1
`define EO3HS_A_R_Z_F 0.1

module EO3HS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   xor  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      if (A && B || !A && !B) (C +=> Z) = (`EO3HS_C_R_Z_R,`EO3HS_C_F_Z_F);
      if (!A && B || A && !B) (C -=> Z) = (`EO3HS_C_F_Z_R,`EO3HS_C_R_Z_F);
      if (A && C || !A && !C) (B +=> Z) = (`EO3HS_B_R_Z_R,`EO3HS_B_F_Z_F);
      if (!A && C || A && !C) (B -=> Z) = (`EO3HS_B_F_Z_R,`EO3HS_B_R_Z_F);
      if (B && C || !B && !C) (A +=> Z) = (`EO3HS_A_R_Z_R,`EO3HS_A_F_Z_F);
      if (!B && C || B && !C) (A -=> Z) = (`EO3HS_A_F_Z_R,`EO3HS_A_R_Z_F);

   endspecify
`endif


endmodule // EO3HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:47 and Version :1.1 //
 
//  START 
// CELL EO3HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define EO3HSP_C_F_Z_F 0.1
`define EO3HSP_C_R_Z_R 0.1
`define EO3HSP_C_F_Z_R 0.1
`define EO3HSP_C_R_Z_F 0.1
`define EO3HSP_B_F_Z_F 0.1
`define EO3HSP_B_R_Z_R 0.1
`define EO3HSP_B_F_Z_R 0.1
`define EO3HSP_B_R_Z_F 0.1
`define EO3HSP_A_F_Z_F 0.1
`define EO3HSP_A_R_Z_R 0.1
`define EO3HSP_A_F_Z_R 0.1
`define EO3HSP_A_R_Z_F 0.1

module EO3HSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   xor  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      if (A && B || !A && !B) (C +=> Z) = (`EO3HSP_C_R_Z_R,`EO3HSP_C_F_Z_F);
      if (!A && B || A && !B) (C -=> Z) = (`EO3HSP_C_F_Z_R,`EO3HSP_C_R_Z_F);
      if (A && C || !A && !C) (B +=> Z) = (`EO3HSP_B_R_Z_R,`EO3HSP_B_F_Z_F);
      if (!A && C || A && !C) (B -=> Z) = (`EO3HSP_B_F_Z_R,`EO3HSP_B_R_Z_F);
      if (B && C || !B && !C) (A +=> Z) = (`EO3HSP_A_R_Z_R,`EO3HSP_A_F_Z_F);
      if (!B && C || B && !C) (A -=> Z) = (`EO3HSP_A_F_Z_R,`EO3HSP_A_R_Z_F);

   endspecify
`endif


endmodule // EO3HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:47 and Version :1.1 //
 
//  START 
// CELL EO3HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define EO3HSX4_C_F_Z_F 0.1
`define EO3HSX4_C_R_Z_R 0.1
`define EO3HSX4_C_F_Z_R 0.1
`define EO3HSX4_C_R_Z_F 0.1
`define EO3HSX4_B_F_Z_F 0.1
`define EO3HSX4_B_R_Z_R 0.1
`define EO3HSX4_B_F_Z_R 0.1
`define EO3HSX4_B_R_Z_F 0.1
`define EO3HSX4_A_F_Z_F 0.1
`define EO3HSX4_A_R_Z_R 0.1
`define EO3HSX4_A_F_Z_R 0.1
`define EO3HSX4_A_R_Z_F 0.1

module EO3HSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   xor  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      if (A && B || !A && !B) (C +=> Z) = (`EO3HSX4_C_R_Z_R,`EO3HSX4_C_F_Z_F);
      if (!A && B || A && !B) (C -=> Z) = (`EO3HSX4_C_F_Z_R,`EO3HSX4_C_R_Z_F);
      if (A && C || !A && !C) (B +=> Z) = (`EO3HSX4_B_R_Z_R,`EO3HSX4_B_F_Z_F);
      if (!A && C || A && !C) (B -=> Z) = (`EO3HSX4_B_F_Z_R,`EO3HSX4_B_R_Z_F);
      if (B && C || !B && !C) (A +=> Z) = (`EO3HSX4_A_R_Z_R,`EO3HSX4_A_F_Z_F);
      if (!B && C || B && !C) (A -=> Z) = (`EO3HSX4_A_F_Z_R,`EO3HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // EO3HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:47 and Version :1.1 //
 
//  START 
// CELL F_EO3HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_EO3HSP_C_F_Z_F 0.1
`define F_EO3HSP_C_R_Z_R 0.1
`define F_EO3HSP_C_F_Z_R 0.1
`define F_EO3HSP_C_R_Z_F 0.1
`define F_EO3HSP_B_F_Z_F 0.1
`define F_EO3HSP_B_R_Z_R 0.1
`define F_EO3HSP_B_F_Z_R 0.1
`define F_EO3HSP_B_R_Z_F 0.1
`define F_EO3HSP_A_F_Z_F 0.1
`define F_EO3HSP_A_R_Z_R 0.1
`define F_EO3HSP_A_F_Z_R 0.1
`define F_EO3HSP_A_R_Z_F 0.1

module F_EO3HSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   xor  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      if (A && B || !A && !B) (C +=> Z) = (`F_EO3HSP_C_R_Z_R,`F_EO3HSP_C_F_Z_F);
      if (!A && B || A && !B) (C -=> Z) = (`F_EO3HSP_C_F_Z_R,`F_EO3HSP_C_R_Z_F);
      if (A && C || !A && !C) (B +=> Z) = (`F_EO3HSP_B_R_Z_R,`F_EO3HSP_B_F_Z_F);
      if (!A && C || A && !C) (B -=> Z) = (`F_EO3HSP_B_F_Z_R,`F_EO3HSP_B_R_Z_F);
      if (B && C || !B && !C) (A +=> Z) = (`F_EO3HSP_A_R_Z_R,`F_EO3HSP_A_F_Z_F);
      if (!B && C || B && !C) (A -=> Z) = (`F_EO3HSP_A_F_Z_R,`F_EO3HSP_A_R_Z_F);

   endspecify
`endif


endmodule // F_EO3HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:47 and Version :1.1 //
 
//  START 
// CELL F_EO3HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_EO3HSX4_C_F_Z_F 0.1
`define F_EO3HSX4_C_R_Z_R 0.1
`define F_EO3HSX4_C_F_Z_R 0.1
`define F_EO3HSX4_C_R_Z_F 0.1
`define F_EO3HSX4_B_F_Z_F 0.1
`define F_EO3HSX4_B_R_Z_R 0.1
`define F_EO3HSX4_B_F_Z_R 0.1
`define F_EO3HSX4_B_R_Z_F 0.1
`define F_EO3HSX4_A_F_Z_F 0.1
`define F_EO3HSX4_A_R_Z_R 0.1
`define F_EO3HSX4_A_F_Z_R 0.1
`define F_EO3HSX4_A_R_Z_F 0.1

module F_EO3HSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   xor  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      if (A && B || !A && !B) (C +=> Z) = (`F_EO3HSX4_C_R_Z_R,`F_EO3HSX4_C_F_Z_F);
      if (!A && B || A && !B) (C -=> Z) = (`F_EO3HSX4_C_F_Z_R,`F_EO3HSX4_C_R_Z_F);
      if (A && C || !A && !C) (B +=> Z) = (`F_EO3HSX4_B_R_Z_R,`F_EO3HSX4_B_F_Z_F);
      if (!A && C || A && !C) (B -=> Z) = (`F_EO3HSX4_B_F_Z_R,`F_EO3HSX4_B_R_Z_F);
      if (B && C || !B && !C) (A +=> Z) = (`F_EO3HSX4_A_R_Z_R,`F_EO3HSX4_A_F_Z_F);
      if (!B && C || B && !C) (A -=> Z) = (`F_EO3HSX4_A_F_Z_R,`F_EO3HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // F_EO3HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:47 and Version :1.1 //
 
//  START 
// CELL FA1HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FA1HS_CI_F_CO_F 0.1
`define FA1HS_CI_R_CO_R 0.1
`define FA1HS_B_F_CO_F 0.1
`define FA1HS_B_R_CO_R 0.1
`define FA1HS_A_F_CO_F 0.1
`define FA1HS_A_R_CO_R 0.1
`define FA1HS_CI_F_Z_F 0.1
`define FA1HS_CI_R_Z_R 0.1
`define FA1HS_CI_F_Z_R 0.1
`define FA1HS_CI_R_Z_F 0.1
`define FA1HS_B_F_Z_F 0.1
`define FA1HS_B_R_Z_R 0.1
`define FA1HS_B_F_Z_R 0.1
`define FA1HS_B_R_Z_F 0.1
`define FA1HS_A_F_Z_F 0.1
`define FA1HS_A_R_Z_R 0.1
`define FA1HS_A_F_Z_R 0.1
`define FA1HS_A_R_Z_F 0.1

module FA1HS (Z, CO, A, B, CI);

   output Z;
   output CO;
   input A;
   input B;
   input CI;


   xor  u0 (Z, A, B, CI);
   // gate-level netlist replaced by UDPs - 19 DEC 1995
   U_MAJ  u1 (CO, A, B, CI);


`ifdef functional
`else
   specify

      (CI +=> CO) = (`FA1HS_CI_R_CO_R,`FA1HS_CI_F_CO_F);
      (B +=> CO) = (`FA1HS_B_R_CO_R,`FA1HS_B_F_CO_F);
      (A +=> CO) = (`FA1HS_A_R_CO_R,`FA1HS_A_F_CO_F);
      if (A && B || !A && !B) (CI +=> Z) = (`FA1HS_CI_R_Z_R,`FA1HS_CI_F_Z_F);
      if (!A && B || A && !B) (CI -=> Z) = (`FA1HS_CI_F_Z_R,`FA1HS_CI_R_Z_F);
      if (A && CI || !A && !CI) (B +=> Z) = (`FA1HS_B_R_Z_R,`FA1HS_B_F_Z_F);
      if (!A && CI || A && !CI) (B -=> Z) = (`FA1HS_B_F_Z_R,`FA1HS_B_R_Z_F);
      if (B && CI || !B && !CI) (A +=> Z) = (`FA1HS_A_R_Z_R,`FA1HS_A_F_Z_F);
      if (!B && CI || B && !CI) (A -=> Z) = (`FA1HS_A_F_Z_R,`FA1HS_A_R_Z_F);

   endspecify
`endif


endmodule // FA1HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:51 and Version :1.1 //
 
//  START 
// CELL FA1HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FA1HSP_CI_F_CO_F 0.1
`define FA1HSP_CI_R_CO_R 0.1
`define FA1HSP_B_F_CO_F 0.1
`define FA1HSP_B_R_CO_R 0.1
`define FA1HSP_A_F_CO_F 0.1
`define FA1HSP_A_R_CO_R 0.1
`define FA1HSP_CI_F_Z_F 0.1
`define FA1HSP_CI_R_Z_R 0.1
`define FA1HSP_CI_F_Z_R 0.1
`define FA1HSP_CI_R_Z_F 0.1
`define FA1HSP_B_F_Z_F 0.1
`define FA1HSP_B_R_Z_R 0.1
`define FA1HSP_B_F_Z_R 0.1
`define FA1HSP_B_R_Z_F 0.1
`define FA1HSP_A_F_Z_F 0.1
`define FA1HSP_A_R_Z_R 0.1
`define FA1HSP_A_F_Z_R 0.1
`define FA1HSP_A_R_Z_F 0.1

module FA1HSP (Z, CO, A, B, CI);

   output Z;
   output CO;
   input A;
   input B;
   input CI;


   xor  u0 (Z, A, B, CI);
   // gate-level netlist replaced by UDPs - 19 DEC 1995
   U_MAJ  u1 (CO, A, B, CI);


`ifdef functional
`else
   specify

      (CI +=> CO) = (`FA1HSP_CI_R_CO_R,`FA1HSP_CI_F_CO_F);
      (B +=> CO) = (`FA1HSP_B_R_CO_R,`FA1HSP_B_F_CO_F);
      (A +=> CO) = (`FA1HSP_A_R_CO_R,`FA1HSP_A_F_CO_F);
      if (A && B || !A && !B) (CI +=> Z) = (`FA1HSP_CI_R_Z_R,`FA1HSP_CI_F_Z_F);
      if (!A && B || A && !B) (CI -=> Z) = (`FA1HSP_CI_F_Z_R,`FA1HSP_CI_R_Z_F);
      if (A && CI || !A && !CI) (B +=> Z) = (`FA1HSP_B_R_Z_R,`FA1HSP_B_F_Z_F);
      if (!A && CI || A && !CI) (B -=> Z) = (`FA1HSP_B_F_Z_R,`FA1HSP_B_R_Z_F);
      if (B && CI || !B && !CI) (A +=> Z) = (`FA1HSP_A_R_Z_R,`FA1HSP_A_F_Z_F);
      if (!B && CI || B && !CI) (A -=> Z) = (`FA1HSP_A_F_Z_R,`FA1HSP_A_R_Z_F);

   endspecify
`endif


endmodule // FA1HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:51 and Version :1.1 //
 
//  START 
// CELL FA1HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FA1HSX4_CI_F_CO_F 0.1
`define FA1HSX4_CI_R_CO_R 0.1
`define FA1HSX4_B_F_CO_F 0.1
`define FA1HSX4_B_R_CO_R 0.1
`define FA1HSX4_A_F_CO_F 0.1
`define FA1HSX4_A_R_CO_R 0.1
`define FA1HSX4_CI_F_Z_F 0.1
`define FA1HSX4_CI_R_Z_R 0.1
`define FA1HSX4_CI_F_Z_R 0.1
`define FA1HSX4_CI_R_Z_F 0.1
`define FA1HSX4_B_F_Z_F 0.1
`define FA1HSX4_B_R_Z_R 0.1
`define FA1HSX4_B_F_Z_R 0.1
`define FA1HSX4_B_R_Z_F 0.1
`define FA1HSX4_A_F_Z_F 0.1
`define FA1HSX4_A_R_Z_R 0.1
`define FA1HSX4_A_F_Z_R 0.1
`define FA1HSX4_A_R_Z_F 0.1

module FA1HSX4 (Z, CO, A, B, CI);

   output Z;
   output CO;
   input A;
   input B;
   input CI;


   xor  u0 (Z, A, B, CI);
   // gate-level netlist replaced by UDPs - 19 DEC 1995
   U_MAJ  u1 (CO, A, B, CI);


`ifdef functional
`else
   specify

      (CI +=> CO) = (`FA1HSX4_CI_R_CO_R,`FA1HSX4_CI_F_CO_F);
      (B +=> CO) = (`FA1HSX4_B_R_CO_R,`FA1HSX4_B_F_CO_F);
      (A +=> CO) = (`FA1HSX4_A_R_CO_R,`FA1HSX4_A_F_CO_F);
      if (A && B || !A && !B) (CI +=> Z) = (`FA1HSX4_CI_R_Z_R,`FA1HSX4_CI_F_Z_F);
      if (!A && B || A && !B) (CI -=> Z) = (`FA1HSX4_CI_F_Z_R,`FA1HSX4_CI_R_Z_F);
      if (A && CI || !A && !CI) (B +=> Z) = (`FA1HSX4_B_R_Z_R,`FA1HSX4_B_F_Z_F);
      if (!A && CI || A && !CI) (B -=> Z) = (`FA1HSX4_B_F_Z_R,`FA1HSX4_B_R_Z_F);
      if (B && CI || !B && !CI) (A +=> Z) = (`FA1HSX4_A_R_Z_R,`FA1HSX4_A_F_Z_F);
      if (!B && CI || B && !CI) (A -=> Z) = (`FA1HSX4_A_F_Z_R,`FA1HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // FA1HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:51 and Version :1.1 //
 
//  START 
// CELL FAS1HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FAS1HSP_CI_F_CO_F 0.1
`define FAS1HSP_CI_R_CO_R 0.1
`define FAS1HSP_B_F_CO_F 0.1
`define FAS1HSP_B_R_CO_R 0.1
`define FAS1HSP_A_F_CO_F 0.1
`define FAS1HSP_A_R_CO_R 0.1
`define FAS1HSP_CI_F_Z_F 0.1
`define FAS1HSP_CI_R_Z_R 0.1
`define FAS1HSP_CI_F_Z_R 0.1
`define FAS1HSP_CI_R_Z_F 0.1
`define FAS1HSP_B_F_Z_F 0.1
`define FAS1HSP_B_R_Z_R 0.1
`define FAS1HSP_B_F_Z_R 0.1
`define FAS1HSP_B_R_Z_F 0.1
`define FAS1HSP_A_F_Z_F 0.1
`define FAS1HSP_A_R_Z_R 0.1
`define FAS1HSP_A_F_Z_R 0.1
`define FAS1HSP_A_R_Z_F 0.1

module FAS1HSP (Z, CO, A, B, CI);

   output Z;
   output CO;
   input A;
   input B;
   input CI;


   xor  u0 (Z, A, B, CI);
   // gate-level netlist replaced by UDPs - 19 DEC 1995
   U_MAJ  u1 (CO, A, B, CI);


`ifdef functional
`else
   specify

      (CI +=> CO) = (`FAS1HSP_CI_R_CO_R,`FAS1HSP_CI_F_CO_F);
      (B +=> CO) = (`FAS1HSP_B_R_CO_R,`FAS1HSP_B_F_CO_F);
      (A +=> CO) = (`FAS1HSP_A_R_CO_R,`FAS1HSP_A_F_CO_F);
      if (A && B || !A && !B) (CI +=> Z) = (`FAS1HSP_CI_R_Z_R,`FAS1HSP_CI_F_Z_F);
      if (!A && B || A && !B) (CI -=> Z) = (`FAS1HSP_CI_F_Z_R,`FAS1HSP_CI_R_Z_F);
      if (A && CI || !A && !CI) (B +=> Z) = (`FAS1HSP_B_R_Z_R,`FAS1HSP_B_F_Z_F);
      if (!A && CI || A && !CI) (B -=> Z) = (`FAS1HSP_B_F_Z_R,`FAS1HSP_B_R_Z_F);
      if (B && CI || !B && !CI) (A +=> Z) = (`FAS1HSP_A_R_Z_R,`FAS1HSP_A_F_Z_F);
      if (!B && CI || B && !CI) (A -=> Z) = (`FAS1HSP_A_F_Z_R,`FAS1HSP_A_R_Z_F);

   endspecify
`endif


endmodule // FAS1HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:51 and Version :1.1 //
 
//  START 
// CELL FAS1HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FAS1HSX4_CI_F_CO_F 0.1
`define FAS1HSX4_CI_R_CO_R 0.1
`define FAS1HSX4_B_F_CO_F 0.1
`define FAS1HSX4_B_R_CO_R 0.1
`define FAS1HSX4_A_F_CO_F 0.1
`define FAS1HSX4_A_R_CO_R 0.1
`define FAS1HSX4_CI_F_Z_F 0.1
`define FAS1HSX4_CI_R_Z_R 0.1
`define FAS1HSX4_CI_F_Z_R 0.1
`define FAS1HSX4_CI_R_Z_F 0.1
`define FAS1HSX4_B_F_Z_F 0.1
`define FAS1HSX4_B_R_Z_R 0.1
`define FAS1HSX4_B_F_Z_R 0.1
`define FAS1HSX4_B_R_Z_F 0.1
`define FAS1HSX4_A_F_Z_F 0.1
`define FAS1HSX4_A_R_Z_R 0.1
`define FAS1HSX4_A_F_Z_R 0.1
`define FAS1HSX4_A_R_Z_F 0.1

module FAS1HSX4 (Z, CO, A, B, CI);

   output Z;
   output CO;
   input A;
   input B;
   input CI;


   xor  u0 (Z, A, B, CI);
   // gate-level netlist replaced by UDPs - 19 DEC 1995
   U_MAJ  u1 (CO, A, B, CI);


`ifdef functional
`else
   specify

      (CI +=> CO) = (`FAS1HSX4_CI_R_CO_R,`FAS1HSX4_CI_F_CO_F);
      (B +=> CO) = (`FAS1HSX4_B_R_CO_R,`FAS1HSX4_B_F_CO_F);
      (A +=> CO) = (`FAS1HSX4_A_R_CO_R,`FAS1HSX4_A_F_CO_F);
      if (A && B || !A && !B) (CI +=> Z) = (`FAS1HSX4_CI_R_Z_R,`FAS1HSX4_CI_F_Z_F);
      if (!A && B || A && !B) (CI -=> Z) = (`FAS1HSX4_CI_F_Z_R,`FAS1HSX4_CI_R_Z_F);
      if (A && CI || !A && !CI) (B +=> Z) = (`FAS1HSX4_B_R_Z_R,`FAS1HSX4_B_F_Z_F);
      if (!A && CI || A && !CI) (B -=> Z) = (`FAS1HSX4_B_F_Z_R,`FAS1HSX4_B_R_Z_F);
      if (B && CI || !B && !CI) (A +=> Z) = (`FAS1HSX4_A_R_Z_R,`FAS1HSX4_A_F_Z_F);
      if (!B && CI || B && !CI) (A -=> Z) = (`FAS1HSX4_A_F_Z_R,`FAS1HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // FAS1HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:51 and Version :1.1 //
 
//  START 
// CELL F_FA1HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_FA1HSP_CI_F_CO_F 0.1
`define F_FA1HSP_CI_R_CO_R 0.1
`define F_FA1HSP_B_F_CO_F 0.1
`define F_FA1HSP_B_R_CO_R 0.1
`define F_FA1HSP_A_F_CO_F 0.1
`define F_FA1HSP_A_R_CO_R 0.1
`define F_FA1HSP_CI_F_Z_F 0.1
`define F_FA1HSP_CI_R_Z_R 0.1
`define F_FA1HSP_CI_F_Z_R 0.1
`define F_FA1HSP_CI_R_Z_F 0.1
`define F_FA1HSP_B_F_Z_F 0.1
`define F_FA1HSP_B_R_Z_R 0.1
`define F_FA1HSP_B_F_Z_R 0.1
`define F_FA1HSP_B_R_Z_F 0.1
`define F_FA1HSP_A_F_Z_F 0.1
`define F_FA1HSP_A_R_Z_R 0.1
`define F_FA1HSP_A_F_Z_R 0.1
`define F_FA1HSP_A_R_Z_F 0.1

module F_FA1HSP (Z, CO, A, B, CI);

   output Z;
   output CO;
   input A;
   input B;
   input CI;


   xor  u0 (Z, A, B, CI);
   // gate-level netlist replaced by UDPs - 19 DEC 1995
   U_MAJ  u1 (CO, A, B, CI);


`ifdef functional
`else
   specify

      (CI +=> CO) = (`F_FA1HSP_CI_R_CO_R,`F_FA1HSP_CI_F_CO_F);
      (B +=> CO) = (`F_FA1HSP_B_R_CO_R,`F_FA1HSP_B_F_CO_F);
      (A +=> CO) = (`F_FA1HSP_A_R_CO_R,`F_FA1HSP_A_F_CO_F);
      if (A && B || !A && !B) (CI +=> Z) = (`F_FA1HSP_CI_R_Z_R,`F_FA1HSP_CI_F_Z_F);
      if (!A && B || A && !B) (CI -=> Z) = (`F_FA1HSP_CI_F_Z_R,`F_FA1HSP_CI_R_Z_F);
      if (A && CI || !A && !CI) (B +=> Z) = (`F_FA1HSP_B_R_Z_R,`F_FA1HSP_B_F_Z_F);
      if (!A && CI || A && !CI) (B -=> Z) = (`F_FA1HSP_B_F_Z_R,`F_FA1HSP_B_R_Z_F);
      if (B && CI || !B && !CI) (A +=> Z) = (`F_FA1HSP_A_R_Z_R,`F_FA1HSP_A_F_Z_F);
      if (!B && CI || B && !CI) (A -=> Z) = (`F_FA1HSP_A_F_Z_R,`F_FA1HSP_A_R_Z_F);

   endspecify
`endif


endmodule // F_FA1HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:51 and Version :1.1 //
 
//  START 
// CELL FA2HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FA2HS_CI_F_CO_F 0.1
`define FA2HS_CI_R_CO_R 0.1
`define FA2HS_B1_F_CO_F 0.1
`define FA2HS_B1_R_CO_R 0.1
`define FA2HS_B0_F_CO_F 0.1
`define FA2HS_B0_R_CO_R 0.1
`define FA2HS_A1_F_CO_F 0.1
`define FA2HS_A1_R_CO_R 0.1
`define FA2HS_A0_F_CO_F 0.1
`define FA2HS_A0_R_CO_R 0.1
`define FA2HS_CI_F_Z1_F 0.1
`define FA2HS_CI_R_Z1_R 0.1
`define FA2HS_CI_F_Z1_R 0.1
`define FA2HS_CI_R_Z1_F 0.1
`define FA2HS_B1_F_Z1_F 0.1
`define FA2HS_B1_R_Z1_R 0.1
`define FA2HS_B1_F_Z1_R 0.1
`define FA2HS_B1_R_Z1_F 0.1
`define FA2HS_B0_F_Z1_F 0.1
`define FA2HS_B0_R_Z1_R 0.1
`define FA2HS_B0_F_Z1_R 0.1
`define FA2HS_B0_R_Z1_F 0.1
`define FA2HS_A1_F_Z1_F 0.1
`define FA2HS_A1_R_Z1_R 0.1
`define FA2HS_A1_F_Z1_R 0.1
`define FA2HS_A1_R_Z1_F 0.1
`define FA2HS_A0_F_Z1_F 0.1
`define FA2HS_A0_R_Z1_R 0.1
`define FA2HS_A0_F_Z1_R 0.1
`define FA2HS_A0_R_Z1_F 0.1
`define FA2HS_CI_F_Z0_F 0.1
`define FA2HS_CI_R_Z0_R 0.1
`define FA2HS_CI_F_Z0_R 0.1
`define FA2HS_CI_R_Z0_F 0.1
`define FA2HS_B0_F_Z0_F 0.1
`define FA2HS_B0_R_Z0_R 0.1
`define FA2HS_B0_F_Z0_R 0.1
`define FA2HS_B0_R_Z0_F 0.1
`define FA2HS_A0_F_Z0_F 0.1
`define FA2HS_A0_R_Z0_R 0.1
`define FA2HS_A0_F_Z0_R 0.1
`define FA2HS_A0_R_Z0_F 0.1

module FA2HS (Z0, Z1, CO, A0, A1, B0, B1, CI);

   output Z0;
   output Z1;
   output CO;
   input A0;
   input A1;
   input B0;
   input B1;
   input CI;


   xor  u0 (Z0, A0, B0, CI);
   xor  u1 (Z1, A1, B1, CO0);
   U_MAJ  u2 (CO, A1, B1, CO0);
   U_MAJ  u3 (CO0, A0, B0, CI);


`ifdef functional
`else
   specify

      (CI +=> CO) = (`FA2HS_CI_R_CO_R,`FA2HS_CI_F_CO_F);
      (B1 +=> CO) = (`FA2HS_B1_R_CO_R,`FA2HS_B1_F_CO_F);
      (B0 +=> CO) = (`FA2HS_B0_R_CO_R,`FA2HS_B0_F_CO_F);
      (A1 +=> CO) = (`FA2HS_A1_R_CO_R,`FA2HS_A1_F_CO_F);
      (A0 +=> CO) = (`FA2HS_A0_R_CO_R,`FA2HS_A0_F_CO_F);
      if (!A0 && A1 && B0 && B1 || A0 && A1 && !B0 && B1 || !A0 && !A1 && B0 && !B1 || A0 && !A1 && !B0 && !B1) (CI +=> Z1) = (`FA2HS_CI_R_Z1_R,`FA2HS_CI_F_Z1_F);
      if (!A0 && !A1 && B0 && B1 || A0 && !A1 && !B0 && B1 || !A0 && A1 && B0 && !B1 || A0 && A1 && !B0 && !B1) (CI -=> Z1) = (`FA2HS_CI_F_Z1_R,`FA2HS_CI_R_Z1_F);
      if (A1 && B0 && CI || A0 && A1 && CI || !A0 && !A1 && !B0 || A0 && A1 && B0 || !A0 && !A1 && !CI || !A1 && !B0 && !CI) (B1 +=> Z1) = (`FA2HS_B1_R_Z1_R,`FA2HS_B1_F_Z1_F);
      if (!A1 && B0 && CI || !A0 && A1 && !B0 || A0 && !A1 && CI || !A0 && A1 && !CI || A0 && !A1 && B0 || A1 && !B0 && !CI) (B1 -=> Z1) = (`FA2HS_B1_F_Z1_R,`FA2HS_B1_R_Z1_F);
      if (!A0 && A1 && B1 && CI || !A0 && !A1 && !B1 && CI || A0 && A1 && B1 && !CI || A0 && !A1 && !B1 && !CI) (B0 +=> Z1) = (`FA2HS_B0_R_Z1_R,`FA2HS_B0_F_Z1_F);
      if (!A0 && !A1 && B1 && CI || !A0 && A1 && !B1 && CI || A0 && !A1 && B1 && !CI || A0 && A1 && !B1 && !CI) (B0 -=> Z1) = (`FA2HS_B0_F_Z1_R,`FA2HS_B0_R_Z1_F);
      if (B0 && B1 && CI || A0 && B1 && CI || !A0 && !B0 && !B1 || A0 && B0 && B1 || !A0 && !B1 && !CI || !B0 && !B1 && !CI) (A1 +=> Z1) = (`FA2HS_A1_R_Z1_R,`FA2HS_A1_F_Z1_F);
      if (!A0 && !B0 && B1 || B0 && !B1 && CI || A0 && !B1 && CI || !A0 && B1 && !CI || !B0 && B1 && !CI || A0 && B0 && !B1) (A1 -=> Z1) = (`FA2HS_A1_F_Z1_R,`FA2HS_A1_R_Z1_F);
      if (A1 && !B0 && B1 && CI || !A1 && !B0 && !B1 && CI || A1 && B0 && B1 && !CI || !A1 && B0 && !B1 && !CI) (A0 +=> Z1) = (`FA2HS_A0_R_Z1_R,`FA2HS_A0_F_Z1_F);
      if (!A1 && !B0 && B1 && CI || A1 && !B0 && !B1 && CI || !A1 && B0 && B1 && !CI || A1 && B0 && !B1 && !CI) (A0 -=> Z1) = (`FA2HS_A0_F_Z1_R,`FA2HS_A0_R_Z1_F);
      if (A0 && B0 || !A0 && !B0) (CI +=> Z0) = (`FA2HS_CI_R_Z0_R,`FA2HS_CI_F_Z0_F);
      if (!A0 && B0 || A0 && !B0) (CI -=> Z0) = (`FA2HS_CI_F_Z0_R,`FA2HS_CI_R_Z0_F);
      if (A0 && CI || !A0 && !CI) (B0 +=> Z0) = (`FA2HS_B0_R_Z0_R,`FA2HS_B0_F_Z0_F);
      if (!A0 && CI || A0 && !CI) (B0 -=> Z0) = (`FA2HS_B0_F_Z0_R,`FA2HS_B0_R_Z0_F);
      if (B0 && CI || !B0 && !CI) (A0 +=> Z0) = (`FA2HS_A0_R_Z0_R,`FA2HS_A0_F_Z0_F);
      if (!B0 && CI || B0 && !CI) (A0 -=> Z0) = (`FA2HS_A0_F_Z0_R,`FA2HS_A0_R_Z0_F);

   endspecify
`endif


endmodule // FA2HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:53 and Version :1.1 //
 
 
//  START 
// CELL FA2HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FA2HSP_CI_F_CO_F 0.1
`define FA2HSP_CI_R_CO_R 0.1
`define FA2HSP_B1_F_CO_F 0.1
`define FA2HSP_B1_R_CO_R 0.1
`define FA2HSP_B0_F_CO_F 0.1
`define FA2HSP_B0_R_CO_R 0.1
`define FA2HSP_A1_F_CO_F 0.1
`define FA2HSP_A1_R_CO_R 0.1
`define FA2HSP_A0_F_CO_F 0.1
`define FA2HSP_A0_R_CO_R 0.1
`define FA2HSP_CI_F_Z1_F 0.1
`define FA2HSP_CI_R_Z1_R 0.1
`define FA2HSP_CI_F_Z1_R 0.1
`define FA2HSP_CI_R_Z1_F 0.1
`define FA2HSP_B1_F_Z1_F 0.1
`define FA2HSP_B1_R_Z1_R 0.1
`define FA2HSP_B1_F_Z1_R 0.1
`define FA2HSP_B1_R_Z1_F 0.1
`define FA2HSP_B0_F_Z1_F 0.1
`define FA2HSP_B0_R_Z1_R 0.1
`define FA2HSP_B0_F_Z1_R 0.1
`define FA2HSP_B0_R_Z1_F 0.1
`define FA2HSP_A1_F_Z1_F 0.1
`define FA2HSP_A1_R_Z1_R 0.1
`define FA2HSP_A1_F_Z1_R 0.1
`define FA2HSP_A1_R_Z1_F 0.1
`define FA2HSP_A0_F_Z1_F 0.1
`define FA2HSP_A0_R_Z1_R 0.1
`define FA2HSP_A0_F_Z1_R 0.1
`define FA2HSP_A0_R_Z1_F 0.1
`define FA2HSP_CI_F_Z0_F 0.1
`define FA2HSP_CI_R_Z0_R 0.1
`define FA2HSP_CI_F_Z0_R 0.1
`define FA2HSP_CI_R_Z0_F 0.1
`define FA2HSP_B0_F_Z0_F 0.1
`define FA2HSP_B0_R_Z0_R 0.1
`define FA2HSP_B0_F_Z0_R 0.1
`define FA2HSP_B0_R_Z0_F 0.1
`define FA2HSP_A0_F_Z0_F 0.1
`define FA2HSP_A0_R_Z0_R 0.1
`define FA2HSP_A0_F_Z0_R 0.1
`define FA2HSP_A0_R_Z0_F 0.1

module FA2HSP (Z0, Z1, CO, A0, A1, B0, B1, CI);

   output Z0;
   output Z1;
   output CO;
   input A0;
   input A1;
   input B0;
   input B1;
   input CI;


   xor  u0 (Z0, A0, B0, CI);
   xor  u1 (Z1, A1, B1, CO0);
   U_MAJ  u2 (CO, A1, B1, CO0);
   U_MAJ  u3 (CO0, A0, B0, CI);


`ifdef functional
`else
   specify

      (CI +=> CO) = (`FA2HSP_CI_R_CO_R,`FA2HSP_CI_F_CO_F);
      (B1 +=> CO) = (`FA2HSP_B1_R_CO_R,`FA2HSP_B1_F_CO_F);
      (B0 +=> CO) = (`FA2HSP_B0_R_CO_R,`FA2HSP_B0_F_CO_F);
      (A1 +=> CO) = (`FA2HSP_A1_R_CO_R,`FA2HSP_A1_F_CO_F);
      (A0 +=> CO) = (`FA2HSP_A0_R_CO_R,`FA2HSP_A0_F_CO_F);
      if (!A0 && A1 && B0 && B1 || A0 && A1 && !B0 && B1 || !A0 && !A1 && B0 && !B1 || A0 && !A1 && !B0 && !B1) (CI +=> Z1) = (`FA2HSP_CI_R_Z1_R,`FA2HSP_CI_F_Z1_F);
      if (!A0 && !A1 && B0 && B1 || A0 && !A1 && !B0 && B1 || !A0 && A1 && B0 && !B1 || A0 && A1 && !B0 && !B1) (CI -=> Z1) = (`FA2HSP_CI_F_Z1_R,`FA2HSP_CI_R_Z1_F);
      if (A1 && B0 && CI || A0 && A1 && CI || !A0 && !A1 && !B0 || A0 && A1 && B0 || !A0 && !A1 && !CI || !A1 && !B0 && !CI) (B1 +=> Z1) = (`FA2HSP_B1_R_Z1_R,`FA2HSP_B1_F_Z1_F);
      if (!A1 && B0 && CI || !A0 && A1 && !B0 || A0 && !A1 && CI || !A0 && A1 && !CI || A0 && !A1 && B0 || A1 && !B0 && !CI) (B1 -=> Z1) = (`FA2HSP_B1_F_Z1_R,`FA2HSP_B1_R_Z1_F);
      if (!A0 && A1 && B1 && CI || !A0 && !A1 && !B1 && CI || A0 && A1 && B1 && !CI || A0 && !A1 && !B1 && !CI) (B0 +=> Z1) = (`FA2HSP_B0_R_Z1_R,`FA2HSP_B0_F_Z1_F);
      if (!A0 && !A1 && B1 && CI || !A0 && A1 && !B1 && CI || A0 && !A1 && B1 && !CI || A0 && A1 && !B1 && !CI) (B0 -=> Z1) = (`FA2HSP_B0_F_Z1_R,`FA2HSP_B0_R_Z1_F);
      if (B0 && B1 && CI || A0 && B1 && CI || !A0 && !B0 && !B1 || A0 && B0 && B1 || !A0 && !B1 && !CI || !B0 && !B1 && !CI) (A1 +=> Z1) = (`FA2HSP_A1_R_Z1_R,`FA2HSP_A1_F_Z1_F);
      if (!A0 && !B0 && B1 || B0 && !B1 && CI || A0 && !B1 && CI || !A0 && B1 && !CI || !B0 && B1 && !CI || A0 && B0 && !B1) (A1 -=> Z1) = (`FA2HSP_A1_F_Z1_R,`FA2HSP_A1_R_Z1_F);
      if (A1 && !B0 && B1 && CI || !A1 && !B0 && !B1 && CI || A1 && B0 && B1 && !CI || !A1 && B0 && !B1 && !CI) (A0 +=> Z1) = (`FA2HSP_A0_R_Z1_R,`FA2HSP_A0_F_Z1_F);
      if (!A1 && !B0 && B1 && CI || A1 && !B0 && !B1 && CI || !A1 && B0 && B1 && !CI || A1 && B0 && !B1 && !CI) (A0 -=> Z1) = (`FA2HSP_A0_F_Z1_R,`FA2HSP_A0_R_Z1_F);
      if (A0 && B0 || !A0 && !B0) (CI +=> Z0) = (`FA2HSP_CI_R_Z0_R,`FA2HSP_CI_F_Z0_F);
      if (!A0 && B0 || A0 && !B0) (CI -=> Z0) = (`FA2HSP_CI_F_Z0_R,`FA2HSP_CI_R_Z0_F);
      if (A0 && CI || !A0 && !CI) (B0 +=> Z0) = (`FA2HSP_B0_R_Z0_R,`FA2HSP_B0_F_Z0_F);
      if (!A0 && CI || A0 && !CI) (B0 -=> Z0) = (`FA2HSP_B0_F_Z0_R,`FA2HSP_B0_R_Z0_F);
      if (B0 && CI || !B0 && !CI) (A0 +=> Z0) = (`FA2HSP_A0_R_Z0_R,`FA2HSP_A0_F_Z0_F);
      if (!B0 && CI || B0 && !CI) (A0 -=> Z0) = (`FA2HSP_A0_F_Z0_R,`FA2HSP_A0_R_Z0_F);

   endspecify
`endif


endmodule // FA2HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:53 and Version :1.1 //
 
 
//  START 
// CELL FD1HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD1HS_CP_R_QN_F 0.1
`define FD1HS_CP_R_QN_R 0.1
`define FD1HS_CP_R_Q_R 0.1
`define FD1HS_CP_R_Q_F 0.1
`define FD1HS_CP_PWH 0.1
`define FD1HS_CP_PWL 0.1
`define FD1HS_D_CP_SETUP_posedge_posedge 0.1
`define FD1HS_D_CP_SETUP_negedge_posedge 0.1
`define FD1HS_D_CP_HOLD_posedge_posedge 0.1
`define FD1HS_D_CP_HOLD_negedge_posedge 0.1

module FD1HS (Q, QN, D, CP);

   output Q;
   output QN;
   input D;
   input CP;


   reg Notifier;


   U_FD_P_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   specify

      (posedge CP => (Q +: D)) = (`FD1HS_CP_R_Q_R, `FD1HS_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`FD1HS_CP_R_QN_R, `FD1HS_CP_R_QN_F);

	$setuphold(posedge CP, posedge D, `FD1HS_D_CP_SETUP_posedge_posedge, `FD1HS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP, negedge D, `FD1HS_D_CP_SETUP_negedge_posedge, `FD1HS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD1HS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1HS_CP_PWH, 0, Notifier);

   endspecify
`endif


endmodule // FD1HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:57 and Version :1.1 //
 
//  START 
// CELL FD1HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD1HSP_CP_R_QN_F 0.1
`define FD1HSP_CP_R_QN_R 0.1
`define FD1HSP_CP_R_Q_R 0.1
`define FD1HSP_CP_R_Q_F 0.1
`define FD1HSP_CP_PWH 0.1
`define FD1HSP_CP_PWL 0.1
`define FD1HSP_D_CP_SETUP_posedge_posedge 0.1
`define FD1HSP_D_CP_SETUP_negedge_posedge 0.1
`define FD1HSP_D_CP_HOLD_posedge_posedge 0.1
`define FD1HSP_D_CP_HOLD_negedge_posedge 0.1

module FD1HSP (Q, QN, D, CP);

   output Q;
   output QN;
   input D;
   input CP;


   reg Notifier;


   U_FD_P_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   specify

      (posedge CP => (Q +: D)) = (`FD1HSP_CP_R_Q_R, `FD1HSP_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`FD1HSP_CP_R_QN_R, `FD1HSP_CP_R_QN_F);

	$setuphold(posedge CP, posedge D, `FD1HSP_D_CP_SETUP_posedge_posedge, `FD1HSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP, negedge D, `FD1HSP_D_CP_SETUP_negedge_posedge, `FD1HSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD1HSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1HSP_CP_PWH, 0, Notifier);

   endspecify
`endif


endmodule // FD1HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:57 and Version :1.1 //
 
//  START 
// CELL FDM1HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDM1HS_CP_R_QN_F 0.1
`define FDM1HS_CP_R_QN_R 0.1
`define FDM1HS_CP_R_Q_R 0.1
`define FDM1HS_CP_R_Q_F 0.1
`define FDM1HS_CP_PWH 0.1
`define FDM1HS_CP_PWL 0.1
`define FDM1HS_D_CP_SETUP_posedge_posedge 0.1
`define FDM1HS_D_CP_SETUP_negedge_posedge 0.1
`define FDM1HS_D_CP_HOLD_posedge_posedge 0.1
`define FDM1HS_D_CP_HOLD_negedge_posedge 0.1

module FDM1HS (Q, QN, D, CP);

   output Q;
   output QN;
   input D;
   input CP;


   reg Notifier;


   U_FD_P_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   specify

      (posedge CP => (Q +: D)) = (`FDM1HS_CP_R_Q_R, `FDM1HS_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`FDM1HS_CP_R_QN_R, `FDM1HS_CP_R_QN_F);

	$setuphold(posedge CP, posedge D, `FDM1HS_D_CP_SETUP_posedge_posedge, `FDM1HS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP, negedge D, `FDM1HS_D_CP_SETUP_negedge_posedge, `FDM1HS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDM1HS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FDM1HS_CP_PWH, 0, Notifier);

   endspecify
`endif


endmodule // FDM1HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:57 and Version :1.1 //
 
//  START 
// CELL FDM1HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDM1HSP_CP_R_QN_F 0.1
`define FDM1HSP_CP_R_QN_R 0.1
`define FDM1HSP_CP_R_Q_R 0.1
`define FDM1HSP_CP_R_Q_F 0.1
`define FDM1HSP_CP_PWH 0.1
`define FDM1HSP_CP_PWL 0.1
`define FDM1HSP_D_CP_SETUP_posedge_posedge 0.1
`define FDM1HSP_D_CP_SETUP_negedge_posedge 0.1
`define FDM1HSP_D_CP_HOLD_posedge_posedge 0.1
`define FDM1HSP_D_CP_HOLD_negedge_posedge 0.1

module FDM1HSP (Q, QN, D, CP);

   output Q;
   output QN;
   input D;
   input CP;


   reg Notifier;


   U_FD_P_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   specify

      (posedge CP => (Q +: D)) = (`FDM1HSP_CP_R_Q_R, `FDM1HSP_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`FDM1HSP_CP_R_QN_R, `FDM1HSP_CP_R_QN_F);

	$setuphold(posedge CP, posedge D, `FDM1HSP_D_CP_SETUP_posedge_posedge, `FDM1HSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP, negedge D, `FDM1HSP_D_CP_SETUP_negedge_posedge, `FDM1HSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDM1HSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FDM1HSP_CP_PWH, 0, Notifier);

   endspecify
`endif


endmodule // FDM1HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:57 and Version :1.1 //
 
//  START 
// CELL F_FD1HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_FD1HS_CP_R_QN_F 0.1
`define F_FD1HS_CP_R_QN_R 0.1
`define F_FD1HS_CP_R_Q_R 0.1
`define F_FD1HS_CP_R_Q_F 0.1
`define F_FD1HS_CP_PWH 0.1
`define F_FD1HS_CP_PWL 0.1
`define F_FD1HS_D_CP_SETUP_posedge_posedge 0.1
`define F_FD1HS_D_CP_SETUP_negedge_posedge 0.1
`define F_FD1HS_D_CP_HOLD_posedge_posedge 0.1
`define F_FD1HS_D_CP_HOLD_negedge_posedge 0.1

module F_FD1HS (Q, QN, D, CP);

   output Q;
   output QN;
   input D;
   input CP;


   reg Notifier;


   U_FD_P_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   specify

      (posedge CP => (Q +: D)) = (`F_FD1HS_CP_R_Q_R, `F_FD1HS_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`F_FD1HS_CP_R_QN_R, `F_FD1HS_CP_R_QN_F);

	$setuphold(posedge CP, posedge D, `F_FD1HS_D_CP_SETUP_posedge_posedge, `F_FD1HS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP, negedge D, `F_FD1HS_D_CP_SETUP_negedge_posedge, `F_FD1HS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `F_FD1HS_CP_PWL, 0, Notifier);
      $width(posedge CP, `F_FD1HS_CP_PWH, 0, Notifier);

   endspecify
`endif


endmodule // F_FD1HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:57 and Version :1.1 //
 
//  START 
// CELL F_FD1HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_FD1HSP_CP_R_QN_F 0.1
`define F_FD1HSP_CP_R_QN_R 0.1
`define F_FD1HSP_CP_R_Q_R 0.1
`define F_FD1HSP_CP_R_Q_F 0.1
`define F_FD1HSP_CP_PWH 0.1
`define F_FD1HSP_CP_PWL 0.1
`define F_FD1HSP_D_CP_SETUP_posedge_posedge 0.1
`define F_FD1HSP_D_CP_SETUP_negedge_posedge 0.1
`define F_FD1HSP_D_CP_HOLD_posedge_posedge 0.1
`define F_FD1HSP_D_CP_HOLD_negedge_posedge 0.1

module F_FD1HSP (Q, QN, D, CP);

   output Q;
   output QN;
   input D;
   input CP;


   reg Notifier;


   U_FD_P_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   specify

      (posedge CP => (Q +: D)) = (`F_FD1HSP_CP_R_Q_R, `F_FD1HSP_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`F_FD1HSP_CP_R_QN_R, `F_FD1HSP_CP_R_QN_F);

	$setuphold(posedge CP, posedge D, `F_FD1HSP_D_CP_SETUP_posedge_posedge, `F_FD1HSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP, negedge D, `F_FD1HSP_D_CP_SETUP_negedge_posedge, `F_FD1HSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `F_FD1HSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `F_FD1HSP_CP_PWH, 0, Notifier);

   endspecify
`endif


endmodule // F_FD1HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:14:57 and Version :1.1 //
 
//  START 
// CELL FD1QHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD1QHS_CP_R_Q_R 0.1
`define FD1QHS_CP_R_Q_F 0.1
`define FD1QHS_CP_PWH 0.1
`define FD1QHS_CP_PWL 0.1
`define FD1QHS_D_CP_SETUP_posedge_posedge 0.1
`define FD1QHS_D_CP_SETUP_negedge_posedge 0.1
`define FD1QHS_D_CP_HOLD_posedge_posedge 0.1
`define FD1QHS_D_CP_HOLD_negedge_posedge 0.1

module FD1QHS (Q, D, CP);

   output Q;
   input D;
   input CP;


   reg Notifier;


   U_FD_P_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify

      (posedge CP => (Q +: D)) = (`FD1QHS_CP_R_Q_R, `FD1QHS_CP_R_Q_F);

	$setuphold(posedge CP, posedge D, `FD1QHS_D_CP_SETUP_posedge_posedge, `FD1QHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP, negedge D, `FD1QHS_D_CP_SETUP_negedge_posedge, `FD1QHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD1QHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1QHS_CP_PWH, 0, Notifier);

   endspecify
`endif


endmodule // FD1QHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:03 and Version :1.1 //
 
//  START 
// CELL FD1QHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD1QHSP_CP_R_Q_R 0.1
`define FD1QHSP_CP_R_Q_F 0.1
`define FD1QHSP_CP_PWH 0.1
`define FD1QHSP_CP_PWL 0.1
`define FD1QHSP_D_CP_SETUP_posedge_posedge 0.1
`define FD1QHSP_D_CP_SETUP_negedge_posedge 0.1
`define FD1QHSP_D_CP_HOLD_posedge_posedge 0.1
`define FD1QHSP_D_CP_HOLD_negedge_posedge 0.1

module FD1QHSP (Q, D, CP);

   output Q;
   input D;
   input CP;


   reg Notifier;


   U_FD_P_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify

      (posedge CP => (Q +: D)) = (`FD1QHSP_CP_R_Q_R, `FD1QHSP_CP_R_Q_F);

	$setuphold(posedge CP, posedge D, `FD1QHSP_D_CP_SETUP_posedge_posedge, `FD1QHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP, negedge D, `FD1QHSP_D_CP_SETUP_negedge_posedge, `FD1QHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD1QHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1QHSP_CP_PWH, 0, Notifier);

   endspecify
`endif


endmodule // FD1QHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:03 and Version :1.1 //
 
//  START 
// CELL FD1QHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD1QHSX4_CP_R_Q_R 0.1
`define FD1QHSX4_CP_R_Q_F 0.1
`define FD1QHSX4_CP_PWH 0.1
`define FD1QHSX4_CP_PWL 0.1
`define FD1QHSX4_D_CP_SETUP_posedge_posedge 0.1
`define FD1QHSX4_D_CP_SETUP_negedge_posedge 0.1
`define FD1QHSX4_D_CP_HOLD_posedge_posedge 0.1
`define FD1QHSX4_D_CP_HOLD_negedge_posedge 0.1

module FD1QHSX4 (Q, D, CP);

   output Q;
   input D;
   input CP;


   reg Notifier;


   U_FD_P_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify

      (posedge CP => (Q +: D)) = (`FD1QHSX4_CP_R_Q_R, `FD1QHSX4_CP_R_Q_F);

	$setuphold(posedge CP, posedge D, `FD1QHSX4_D_CP_SETUP_posedge_posedge, `FD1QHSX4_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP, negedge D, `FD1QHSX4_D_CP_SETUP_negedge_posedge, `FD1QHSX4_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD1QHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1QHSX4_CP_PWH, 0, Notifier);

   endspecify
`endif


endmodule // FD1QHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:03 and Version :1.1 //
 
//  START 
// CELL FDM1QHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDM1QHS_CP_R_Q_R 0.1
`define FDM1QHS_CP_R_Q_F 0.1
`define FDM1QHS_CP_PWH 0.1
`define FDM1QHS_CP_PWL 0.1
`define FDM1QHS_D_CP_SETUP_posedge_posedge 0.1
`define FDM1QHS_D_CP_SETUP_negedge_posedge 0.1
`define FDM1QHS_D_CP_HOLD_posedge_posedge 0.1
`define FDM1QHS_D_CP_HOLD_negedge_posedge 0.1

module FDM1QHS (Q, D, CP);

   output Q;
   input D;
   input CP;


   reg Notifier;


   U_FD_P_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify

      (posedge CP => (Q +: D)) = (`FDM1QHS_CP_R_Q_R, `FDM1QHS_CP_R_Q_F);

	$setuphold(posedge CP, posedge D, `FDM1QHS_D_CP_SETUP_posedge_posedge, `FDM1QHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP, negedge D, `FDM1QHS_D_CP_SETUP_negedge_posedge, `FDM1QHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDM1QHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FDM1QHS_CP_PWH, 0, Notifier);

   endspecify
`endif


endmodule // FDM1QHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:03 and Version :1.1 //
 
//  START 
// CELL FDM1QHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDM1QHSP_CP_R_Q_R 0.1
`define FDM1QHSP_CP_R_Q_F 0.1
`define FDM1QHSP_CP_PWH 0.1
`define FDM1QHSP_CP_PWL 0.1
`define FDM1QHSP_D_CP_SETUP_posedge_posedge 0.1
`define FDM1QHSP_D_CP_SETUP_negedge_posedge 0.1
`define FDM1QHSP_D_CP_HOLD_posedge_posedge 0.1
`define FDM1QHSP_D_CP_HOLD_negedge_posedge 0.1

module FDM1QHSP (Q, D, CP);

   output Q;
   input D;
   input CP;


   reg Notifier;


   U_FD_P_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify

      (posedge CP => (Q +: D)) = (`FDM1QHSP_CP_R_Q_R, `FDM1QHSP_CP_R_Q_F);

	$setuphold(posedge CP, posedge D, `FDM1QHSP_D_CP_SETUP_posedge_posedge, `FDM1QHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP, negedge D, `FDM1QHSP_D_CP_SETUP_negedge_posedge, `FDM1QHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDM1QHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FDM1QHSP_CP_PWH, 0, Notifier);

   endspecify
`endif


endmodule // FDM1QHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:03 and Version :1.1 //
 
//  START 
// CELL F_FD1QHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_FD1QHS_CP_R_Q_R 0.1
`define F_FD1QHS_CP_R_Q_F 0.1
`define F_FD1QHS_CP_PWH 0.1
`define F_FD1QHS_CP_PWL 0.1
`define F_FD1QHS_D_CP_SETUP_posedge_posedge 0.1
`define F_FD1QHS_D_CP_SETUP_negedge_posedge 0.1
`define F_FD1QHS_D_CP_HOLD_posedge_posedge 0.1
`define F_FD1QHS_D_CP_HOLD_negedge_posedge 0.1

module F_FD1QHS (Q, D, CP);

   output Q;
   input D;
   input CP;


   reg Notifier;


   U_FD_P_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify

      (posedge CP => (Q +: D)) = (`F_FD1QHS_CP_R_Q_R, `F_FD1QHS_CP_R_Q_F);

	$setuphold(posedge CP, posedge D, `F_FD1QHS_D_CP_SETUP_posedge_posedge, `F_FD1QHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP, negedge D, `F_FD1QHS_D_CP_SETUP_negedge_posedge, `F_FD1QHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `F_FD1QHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `F_FD1QHS_CP_PWH, 0, Notifier);

   endspecify
`endif


endmodule // F_FD1QHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:03 and Version :1.1 //
 
//  START 
// CELL F_FD1QHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_FD1QHSP_CP_R_Q_R 0.1
`define F_FD1QHSP_CP_R_Q_F 0.1
`define F_FD1QHSP_CP_PWH 0.1
`define F_FD1QHSP_CP_PWL 0.1
`define F_FD1QHSP_D_CP_SETUP_posedge_posedge 0.1
`define F_FD1QHSP_D_CP_SETUP_negedge_posedge 0.1
`define F_FD1QHSP_D_CP_HOLD_posedge_posedge 0.1
`define F_FD1QHSP_D_CP_HOLD_negedge_posedge 0.1

module F_FD1QHSP (Q, D, CP);

   output Q;
   input D;
   input CP;


   reg Notifier;


   U_FD_P_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify

      (posedge CP => (Q +: D)) = (`F_FD1QHSP_CP_R_Q_R, `F_FD1QHSP_CP_R_Q_F);

	$setuphold(posedge CP, posedge D, `F_FD1QHSP_D_CP_SETUP_posedge_posedge, `F_FD1QHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP, negedge D, `F_FD1QHSP_D_CP_SETUP_negedge_posedge, `F_FD1QHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `F_FD1QHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `F_FD1QHSP_CP_PWH, 0, Notifier);

   endspecify
`endif


endmodule // F_FD1QHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:03 and Version :1.1 //
 
//  START 
// CELL F_FD1QHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_FD1QHSX4_CP_R_Q_R 0.1
`define F_FD1QHSX4_CP_R_Q_F 0.1
`define F_FD1QHSX4_CP_PWH 0.1
`define F_FD1QHSX4_CP_PWL 0.1
`define F_FD1QHSX4_D_CP_SETUP_posedge_posedge 0.1
`define F_FD1QHSX4_D_CP_SETUP_negedge_posedge 0.1
`define F_FD1QHSX4_D_CP_HOLD_posedge_posedge 0.1
`define F_FD1QHSX4_D_CP_HOLD_negedge_posedge 0.1

module F_FD1QHSX4 (Q, D, CP);

   output Q;
   input D;
   input CP;


   reg Notifier;


   U_FD_P_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify

      (posedge CP => (Q +: D)) = (`F_FD1QHSX4_CP_R_Q_R, `F_FD1QHSX4_CP_R_Q_F);

	$setuphold(posedge CP, posedge D, `F_FD1QHSX4_D_CP_SETUP_posedge_posedge, `F_FD1QHSX4_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP, negedge D, `F_FD1QHSX4_D_CP_SETUP_negedge_posedge, `F_FD1QHSX4_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `F_FD1QHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP, `F_FD1QHSX4_CP_PWH, 0, Notifier);

   endspecify
`endif


endmodule // F_FD1QHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:03 and Version :1.1 //
 
//  START 
// CELL FD1SHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD1SHS_CP_R_QN_F 0.1
`define FD1SHS_CP_R_QN_R 0.1
`define FD1SHS_CP_R_Q_R 0.1
`define FD1SHS_CP_R_Q_F 0.1
`define FD1SHS_CP_PWH 0.1
`define FD1SHS_CP_PWL 0.1
`define FD1SHS_D_CP_SETUP_posedge_posedge 0.1
`define FD1SHS_D_CP_SETUP_negedge_posedge 0.1
`define FD1SHS_D_CP_HOLD_posedge_posedge 0.1
`define FD1SHS_D_CP_HOLD_negedge_posedge 0.1
`define FD1SHS_TI_CP_SETUP_posedge_posedge 0.1
`define FD1SHS_TI_CP_SETUP_negedge_posedge 0.1
`define FD1SHS_TI_CP_HOLD_posedge_posedge 0.1
`define FD1SHS_TI_CP_HOLD_negedge_posedge 0.1
`define FD1SHS_TE_CP_SETUP_posedge_posedge 0.1
`define FD1SHS_TE_CP_SETUP_negedge_posedge 0.1
`define FD1SHS_TE_CP_HOLD_posedge_posedge 0.1
`define FD1SHS_TE_CP_HOLD_negedge_posedge 0.1

module FD1SHS (Q, QN, D, CP, TI, TE);

   output Q;
   output QN;
   input D;
   input CP;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault

      if(!TE) (posedge CP => (Q +: D)) = (`FD1SHS_CP_R_Q_R, `FD1SHS_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD1SHS_CP_R_Q_R, `FD1SHS_CP_R_Q_F);
      if(!D && TI) (posedge CP => (Q +: TE)) = (`FD1SHS_CP_R_Q_R, `FD1SHS_CP_R_Q_F);
      if(!TI && D) (posedge CP => (Q -: TE)) = (`FD1SHS_CP_R_Q_R, `FD1SHS_CP_R_Q_F);
      if(!TE) (posedge CP => (QN -: D)) = (`FD1SHS_CP_R_QN_R, `FD1SHS_CP_R_QN_F);
      if(TE) (posedge CP => (QN -: TI)) = (`FD1SHS_CP_R_QN_R, `FD1SHS_CP_R_QN_F);
      if(!D && TI) (posedge CP => (QN -: TE)) = (`FD1SHS_CP_R_QN_R, `FD1SHS_CP_R_QN_F);
      if(!TI && D) (posedge CP => (QN +: TE)) = (`FD1SHS_CP_R_QN_R, `FD1SHS_CP_R_QN_F);

	$setuphold(posedge CP &&& XorDTI_, posedge TE, `FD1SHS_TE_CP_SETUP_posedge_posedge, `FD1SHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& XorDTI_, negedge TE, `FD1SHS_TE_CP_SETUP_negedge_posedge, `FD1SHS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FD1SHS_TI_CP_SETUP_posedge_posedge, `FD1SHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FD1SHS_TI_CP_SETUP_negedge_posedge, `FD1SHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TEX, posedge D, `FD1SHS_D_CP_SETUP_posedge_posedge, `FD1SHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TEX, negedge D, `FD1SHS_D_CP_SETUP_negedge_posedge, `FD1SHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD1SHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1SHS_CP_PWH, 0, Notifier);
`else
     (posedge CP => (Q +: Mux21DTITE_)) = (`FD1SHS_CP_R_Q_R, `FD1SHS_CP_R_Q_F);
     (posedge CP => (QN -: Mux21DTITE_)) = (`FD1SHS_CP_R_QN_R, `FD1SHS_CP_R_QN_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `FD1SHS_TE_CP_SETUP_posedge_posedge, `FD1SHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `FD1SHS_TE_CP_SETUP_negedge_posedge, `FD1SHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD1SHS_TI_CP_SETUP_posedge_posedge, `FD1SHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD1SHS_TI_CP_SETUP_negedge_posedge, `FD1SHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `FD1SHS_D_CP_SETUP_posedge_posedge, `FD1SHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `FD1SHS_D_CP_SETUP_negedge_posedge, `FD1SHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD1SHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1SHS_CP_PWH, 0, Notifier);
`endif 
   endspecify
`endif


endmodule // FD1SHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:07 and Version :1.1 //
 
//  START 

// CELL FD1SHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD1SHSP_CP_R_QN_F 0.1
`define FD1SHSP_CP_R_QN_R 0.1
`define FD1SHSP_CP_R_Q_R 0.1
`define FD1SHSP_CP_R_Q_F 0.1
`define FD1SHSP_CP_PWH 0.1
`define FD1SHSP_CP_PWL 0.1
`define FD1SHSP_D_CP_SETUP_posedge_posedge 0.1
`define FD1SHSP_D_CP_SETUP_negedge_posedge 0.1
`define FD1SHSP_D_CP_HOLD_posedge_posedge 0.1
`define FD1SHSP_D_CP_HOLD_negedge_posedge 0.1
`define FD1SHSP_TI_CP_SETUP_posedge_posedge 0.1
`define FD1SHSP_TI_CP_SETUP_negedge_posedge 0.1
`define FD1SHSP_TI_CP_HOLD_posedge_posedge 0.1
`define FD1SHSP_TI_CP_HOLD_negedge_posedge 0.1
`define FD1SHSP_TE_CP_SETUP_posedge_posedge 0.1
`define FD1SHSP_TE_CP_SETUP_negedge_posedge 0.1
`define FD1SHSP_TE_CP_HOLD_posedge_posedge 0.1
`define FD1SHSP_TE_CP_HOLD_negedge_posedge 0.1

module FD1SHSP (Q, QN, D, CP, TI, TE);

   output Q;
   output QN;
   input D;
   input CP;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault

      if(!TE) (posedge CP => (Q +: D)) = (`FD1SHSP_CP_R_Q_R, `FD1SHSP_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD1SHSP_CP_R_Q_R, `FD1SHSP_CP_R_Q_F);
      if(!D && TI) (posedge CP => (Q +: TE)) = (`FD1SHSP_CP_R_Q_R, `FD1SHSP_CP_R_Q_F);
      if(!TI && D) (posedge CP => (Q -: TE)) = (`FD1SHSP_CP_R_Q_R, `FD1SHSP_CP_R_Q_F);
      if(!TE) (posedge CP => (QN -: D)) = (`FD1SHSP_CP_R_QN_R, `FD1SHSP_CP_R_QN_F);
      if(TE) (posedge CP => (QN -: TI)) = (`FD1SHSP_CP_R_QN_R, `FD1SHSP_CP_R_QN_F);
      if(!D && TI) (posedge CP => (QN -: TE)) = (`FD1SHSP_CP_R_QN_R, `FD1SHSP_CP_R_QN_F);
      if(!TI && D) (posedge CP => (QN +: TE)) = (`FD1SHSP_CP_R_QN_R, `FD1SHSP_CP_R_QN_F);

	$setuphold(posedge CP &&& XorDTI_, posedge TE, `FD1SHSP_TE_CP_SETUP_posedge_posedge, `FD1SHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& XorDTI_, negedge TE, `FD1SHSP_TE_CP_SETUP_negedge_posedge, `FD1SHSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FD1SHSP_TI_CP_SETUP_posedge_posedge, `FD1SHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FD1SHSP_TI_CP_SETUP_negedge_posedge, `FD1SHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TEX, posedge D, `FD1SHSP_D_CP_SETUP_posedge_posedge, `FD1SHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TEX, negedge D, `FD1SHSP_D_CP_SETUP_negedge_posedge, `FD1SHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD1SHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1SHSP_CP_PWH, 0, Notifier);
`else
     (posedge CP => (Q +: Mux21DTITE_)) = (`FD1SHSP_CP_R_Q_R, `FD1SHSP_CP_R_Q_F);
     (posedge CP => (QN -: Mux21DTITE_)) = (`FD1SHSP_CP_R_QN_R, `FD1SHSP_CP_R_QN_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `FD1SHSP_TE_CP_SETUP_posedge_posedge, `FD1SHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `FD1SHSP_TE_CP_SETUP_negedge_posedge, `FD1SHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD1SHSP_TI_CP_SETUP_posedge_posedge, `FD1SHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD1SHSP_TI_CP_SETUP_negedge_posedge, `FD1SHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `FD1SHSP_D_CP_SETUP_posedge_posedge, `FD1SHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `FD1SHSP_D_CP_SETUP_negedge_posedge, `FD1SHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD1SHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1SHSP_CP_PWH, 0, Notifier);
`endif 
   endspecify
`endif


endmodule // FD1SHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:07 and Version :1.1 //
 
//  START 

// CELL FDM1SHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDM1SHS_CP_R_QN_F 0.1
`define FDM1SHS_CP_R_QN_R 0.1
`define FDM1SHS_CP_R_Q_R 0.1
`define FDM1SHS_CP_R_Q_F 0.1
`define FDM1SHS_CP_PWH 0.1
`define FDM1SHS_CP_PWL 0.1
`define FDM1SHS_D_CP_SETUP_posedge_posedge 0.1
`define FDM1SHS_D_CP_SETUP_negedge_posedge 0.1
`define FDM1SHS_D_CP_HOLD_posedge_posedge 0.1
`define FDM1SHS_D_CP_HOLD_negedge_posedge 0.1
`define FDM1SHS_TI_CP_SETUP_posedge_posedge 0.1
`define FDM1SHS_TI_CP_SETUP_negedge_posedge 0.1
`define FDM1SHS_TI_CP_HOLD_posedge_posedge 0.1
`define FDM1SHS_TI_CP_HOLD_negedge_posedge 0.1
`define FDM1SHS_TE_CP_SETUP_posedge_posedge 0.1
`define FDM1SHS_TE_CP_SETUP_negedge_posedge 0.1
`define FDM1SHS_TE_CP_HOLD_posedge_posedge 0.1
`define FDM1SHS_TE_CP_HOLD_negedge_posedge 0.1

module FDM1SHS (Q, QN, D, CP, TI, TE);

   output Q;
   output QN;
   input D;
   input CP;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault

      if(!TE) (posedge CP => (Q +: D)) = (`FDM1SHS_CP_R_Q_R, `FDM1SHS_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FDM1SHS_CP_R_Q_R, `FDM1SHS_CP_R_Q_F);
      if(!D && TI) (posedge CP => (Q +: TE)) = (`FDM1SHS_CP_R_Q_R, `FDM1SHS_CP_R_Q_F);
      if(!TI && D) (posedge CP => (Q -: TE)) = (`FDM1SHS_CP_R_Q_R, `FDM1SHS_CP_R_Q_F);
      if(!TE) (posedge CP => (QN -: D)) = (`FDM1SHS_CP_R_QN_R, `FDM1SHS_CP_R_QN_F);
      if(TE) (posedge CP => (QN -: TI)) = (`FDM1SHS_CP_R_QN_R, `FDM1SHS_CP_R_QN_F);
      if(!D && TI) (posedge CP => (QN -: TE)) = (`FDM1SHS_CP_R_QN_R, `FDM1SHS_CP_R_QN_F);
      if(!TI && D) (posedge CP => (QN +: TE)) = (`FDM1SHS_CP_R_QN_R, `FDM1SHS_CP_R_QN_F);

	$setuphold(posedge CP &&& XorDTI_, posedge TE, `FDM1SHS_TE_CP_SETUP_posedge_posedge, `FDM1SHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& XorDTI_, negedge TE, `FDM1SHS_TE_CP_SETUP_negedge_posedge, `FDM1SHS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FDM1SHS_TI_CP_SETUP_posedge_posedge, `FDM1SHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FDM1SHS_TI_CP_SETUP_negedge_posedge, `FDM1SHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TEX, posedge D, `FDM1SHS_D_CP_SETUP_posedge_posedge, `FDM1SHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TEX, negedge D, `FDM1SHS_D_CP_SETUP_negedge_posedge, `FDM1SHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDM1SHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FDM1SHS_CP_PWH, 0, Notifier);
`else
     (posedge CP => (Q +: Mux21DTITE_)) = (`FDM1SHS_CP_R_Q_R, `FDM1SHS_CP_R_Q_F);
     (posedge CP => (QN -: Mux21DTITE_)) = (`FDM1SHS_CP_R_QN_R, `FDM1SHS_CP_R_QN_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `FDM1SHS_TE_CP_SETUP_posedge_posedge, `FDM1SHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `FDM1SHS_TE_CP_SETUP_negedge_posedge, `FDM1SHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FDM1SHS_TI_CP_SETUP_posedge_posedge, `FDM1SHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FDM1SHS_TI_CP_SETUP_negedge_posedge, `FDM1SHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `FDM1SHS_D_CP_SETUP_posedge_posedge, `FDM1SHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `FDM1SHS_D_CP_SETUP_negedge_posedge, `FDM1SHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDM1SHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FDM1SHS_CP_PWH, 0, Notifier);
`endif 
   endspecify
`endif


endmodule // FDM1SHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:07 and Version :1.1 //
 
//  START 

// CELL FDM1SHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDM1SHSP_CP_R_QN_F 0.1
`define FDM1SHSP_CP_R_QN_R 0.1
`define FDM1SHSP_CP_R_Q_R 0.1
`define FDM1SHSP_CP_R_Q_F 0.1
`define FDM1SHSP_CP_PWH 0.1
`define FDM1SHSP_CP_PWL 0.1
`define FDM1SHSP_D_CP_SETUP_posedge_posedge 0.1
`define FDM1SHSP_D_CP_SETUP_negedge_posedge 0.1
`define FDM1SHSP_D_CP_HOLD_posedge_posedge 0.1
`define FDM1SHSP_D_CP_HOLD_negedge_posedge 0.1
`define FDM1SHSP_TI_CP_SETUP_posedge_posedge 0.1
`define FDM1SHSP_TI_CP_SETUP_negedge_posedge 0.1
`define FDM1SHSP_TI_CP_HOLD_posedge_posedge 0.1
`define FDM1SHSP_TI_CP_HOLD_negedge_posedge 0.1
`define FDM1SHSP_TE_CP_SETUP_posedge_posedge 0.1
`define FDM1SHSP_TE_CP_SETUP_negedge_posedge 0.1
`define FDM1SHSP_TE_CP_HOLD_posedge_posedge 0.1
`define FDM1SHSP_TE_CP_HOLD_negedge_posedge 0.1

module FDM1SHSP (Q, QN, D, CP, TI, TE);

   output Q;
   output QN;
   input D;
   input CP;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault

      if(!TE) (posedge CP => (Q +: D)) = (`FDM1SHSP_CP_R_Q_R, `FDM1SHSP_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FDM1SHSP_CP_R_Q_R, `FDM1SHSP_CP_R_Q_F);
      if(!D && TI) (posedge CP => (Q +: TE)) = (`FDM1SHSP_CP_R_Q_R, `FDM1SHSP_CP_R_Q_F);
      if(!TI && D) (posedge CP => (Q -: TE)) = (`FDM1SHSP_CP_R_Q_R, `FDM1SHSP_CP_R_Q_F);
      if(!TE) (posedge CP => (QN -: D)) = (`FDM1SHSP_CP_R_QN_R, `FDM1SHSP_CP_R_QN_F);
      if(TE) (posedge CP => (QN -: TI)) = (`FDM1SHSP_CP_R_QN_R, `FDM1SHSP_CP_R_QN_F);
      if(!D && TI) (posedge CP => (QN -: TE)) = (`FDM1SHSP_CP_R_QN_R, `FDM1SHSP_CP_R_QN_F);
      if(!TI && D) (posedge CP => (QN +: TE)) = (`FDM1SHSP_CP_R_QN_R, `FDM1SHSP_CP_R_QN_F);

	$setuphold(posedge CP &&& XorDTI_, posedge TE, `FDM1SHSP_TE_CP_SETUP_posedge_posedge, `FDM1SHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& XorDTI_, negedge TE, `FDM1SHSP_TE_CP_SETUP_negedge_posedge, `FDM1SHSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FDM1SHSP_TI_CP_SETUP_posedge_posedge, `FDM1SHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FDM1SHSP_TI_CP_SETUP_negedge_posedge, `FDM1SHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TEX, posedge D, `FDM1SHSP_D_CP_SETUP_posedge_posedge, `FDM1SHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TEX, negedge D, `FDM1SHSP_D_CP_SETUP_negedge_posedge, `FDM1SHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDM1SHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FDM1SHSP_CP_PWH, 0, Notifier);
`else
     (posedge CP => (Q +: Mux21DTITE_)) = (`FDM1SHSP_CP_R_Q_R, `FDM1SHSP_CP_R_Q_F);
     (posedge CP => (QN -: Mux21DTITE_)) = (`FDM1SHSP_CP_R_QN_R, `FDM1SHSP_CP_R_QN_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `FDM1SHSP_TE_CP_SETUP_posedge_posedge, `FDM1SHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `FDM1SHSP_TE_CP_SETUP_negedge_posedge, `FDM1SHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FDM1SHSP_TI_CP_SETUP_posedge_posedge, `FDM1SHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FDM1SHSP_TI_CP_SETUP_negedge_posedge, `FDM1SHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `FDM1SHSP_D_CP_SETUP_posedge_posedge, `FDM1SHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `FDM1SHSP_D_CP_SETUP_negedge_posedge, `FDM1SHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDM1SHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FDM1SHSP_CP_PWH, 0, Notifier);
`endif 
   endspecify
`endif


endmodule // FDM1SHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:07 and Version :1.1 //
 
//  START 

// CELL F_FD1SHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_FD1SHS_CP_R_QN_F 0.1
`define F_FD1SHS_CP_R_QN_R 0.1
`define F_FD1SHS_CP_R_Q_R 0.1
`define F_FD1SHS_CP_R_Q_F 0.1
`define F_FD1SHS_CP_PWH 0.1
`define F_FD1SHS_CP_PWL 0.1
`define F_FD1SHS_D_CP_SETUP_posedge_posedge 0.1
`define F_FD1SHS_D_CP_SETUP_negedge_posedge 0.1
`define F_FD1SHS_D_CP_HOLD_posedge_posedge 0.1
`define F_FD1SHS_D_CP_HOLD_negedge_posedge 0.1
`define F_FD1SHS_TI_CP_SETUP_posedge_posedge 0.1
`define F_FD1SHS_TI_CP_SETUP_negedge_posedge 0.1
`define F_FD1SHS_TI_CP_HOLD_posedge_posedge 0.1
`define F_FD1SHS_TI_CP_HOLD_negedge_posedge 0.1
`define F_FD1SHS_TE_CP_SETUP_posedge_posedge 0.1
`define F_FD1SHS_TE_CP_SETUP_negedge_posedge 0.1
`define F_FD1SHS_TE_CP_HOLD_posedge_posedge 0.1
`define F_FD1SHS_TE_CP_HOLD_negedge_posedge 0.1

module F_FD1SHS (Q, QN, D, CP, TI, TE);

   output Q;
   output QN;
   input D;
   input CP;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault

      if(!TE) (posedge CP => (Q +: D)) = (`F_FD1SHS_CP_R_Q_R, `F_FD1SHS_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`F_FD1SHS_CP_R_Q_R, `F_FD1SHS_CP_R_Q_F);
      if(!D && TI) (posedge CP => (Q +: TE)) = (`F_FD1SHS_CP_R_Q_R, `F_FD1SHS_CP_R_Q_F);
      if(!TI && D) (posedge CP => (Q -: TE)) = (`F_FD1SHS_CP_R_Q_R, `F_FD1SHS_CP_R_Q_F);
      if(!TE) (posedge CP => (QN -: D)) = (`F_FD1SHS_CP_R_QN_R, `F_FD1SHS_CP_R_QN_F);
      if(TE) (posedge CP => (QN -: TI)) = (`F_FD1SHS_CP_R_QN_R, `F_FD1SHS_CP_R_QN_F);
      if(!D && TI) (posedge CP => (QN -: TE)) = (`F_FD1SHS_CP_R_QN_R, `F_FD1SHS_CP_R_QN_F);
      if(!TI && D) (posedge CP => (QN +: TE)) = (`F_FD1SHS_CP_R_QN_R, `F_FD1SHS_CP_R_QN_F);

	$setuphold(posedge CP &&& XorDTI_, posedge TE, `F_FD1SHS_TE_CP_SETUP_posedge_posedge, `F_FD1SHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& XorDTI_, negedge TE, `F_FD1SHS_TE_CP_SETUP_negedge_posedge, `F_FD1SHS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `F_FD1SHS_TI_CP_SETUP_posedge_posedge, `F_FD1SHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `F_FD1SHS_TI_CP_SETUP_negedge_posedge, `F_FD1SHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TEX, posedge D, `F_FD1SHS_D_CP_SETUP_posedge_posedge, `F_FD1SHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TEX, negedge D, `F_FD1SHS_D_CP_SETUP_negedge_posedge, `F_FD1SHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `F_FD1SHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `F_FD1SHS_CP_PWH, 0, Notifier);
`else
     (posedge CP => (Q +: Mux21DTITE_)) = (`F_FD1SHS_CP_R_Q_R, `F_FD1SHS_CP_R_Q_F);
     (posedge CP => (QN -: Mux21DTITE_)) = (`F_FD1SHS_CP_R_QN_R, `F_FD1SHS_CP_R_QN_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `F_FD1SHS_TE_CP_SETUP_posedge_posedge, `F_FD1SHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `F_FD1SHS_TE_CP_SETUP_negedge_posedge, `F_FD1SHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `F_FD1SHS_TI_CP_SETUP_posedge_posedge, `F_FD1SHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `F_FD1SHS_TI_CP_SETUP_negedge_posedge, `F_FD1SHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `F_FD1SHS_D_CP_SETUP_posedge_posedge, `F_FD1SHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `F_FD1SHS_D_CP_SETUP_negedge_posedge, `F_FD1SHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `F_FD1SHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `F_FD1SHS_CP_PWH, 0, Notifier);
`endif 
   endspecify
`endif


endmodule // F_FD1SHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:07 and Version :1.1 //
 
//  START 

// CELL F_FD1SHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_FD1SHSP_CP_R_QN_F 0.1
`define F_FD1SHSP_CP_R_QN_R 0.1
`define F_FD1SHSP_CP_R_Q_R 0.1
`define F_FD1SHSP_CP_R_Q_F 0.1
`define F_FD1SHSP_CP_PWH 0.1
`define F_FD1SHSP_CP_PWL 0.1
`define F_FD1SHSP_D_CP_SETUP_posedge_posedge 0.1
`define F_FD1SHSP_D_CP_SETUP_negedge_posedge 0.1
`define F_FD1SHSP_D_CP_HOLD_posedge_posedge 0.1
`define F_FD1SHSP_D_CP_HOLD_negedge_posedge 0.1
`define F_FD1SHSP_TI_CP_SETUP_posedge_posedge 0.1
`define F_FD1SHSP_TI_CP_SETUP_negedge_posedge 0.1
`define F_FD1SHSP_TI_CP_HOLD_posedge_posedge 0.1
`define F_FD1SHSP_TI_CP_HOLD_negedge_posedge 0.1
`define F_FD1SHSP_TE_CP_SETUP_posedge_posedge 0.1
`define F_FD1SHSP_TE_CP_SETUP_negedge_posedge 0.1
`define F_FD1SHSP_TE_CP_HOLD_posedge_posedge 0.1
`define F_FD1SHSP_TE_CP_HOLD_negedge_posedge 0.1

module F_FD1SHSP (Q, QN, D, CP, TI, TE);

   output Q;
   output QN;
   input D;
   input CP;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault

      if(!TE) (posedge CP => (Q +: D)) = (`F_FD1SHSP_CP_R_Q_R, `F_FD1SHSP_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`F_FD1SHSP_CP_R_Q_R, `F_FD1SHSP_CP_R_Q_F);
      if(!D && TI) (posedge CP => (Q +: TE)) = (`F_FD1SHSP_CP_R_Q_R, `F_FD1SHSP_CP_R_Q_F);
      if(!TI && D) (posedge CP => (Q -: TE)) = (`F_FD1SHSP_CP_R_Q_R, `F_FD1SHSP_CP_R_Q_F);
      if(!TE) (posedge CP => (QN -: D)) = (`F_FD1SHSP_CP_R_QN_R, `F_FD1SHSP_CP_R_QN_F);
      if(TE) (posedge CP => (QN -: TI)) = (`F_FD1SHSP_CP_R_QN_R, `F_FD1SHSP_CP_R_QN_F);
      if(!D && TI) (posedge CP => (QN -: TE)) = (`F_FD1SHSP_CP_R_QN_R, `F_FD1SHSP_CP_R_QN_F);
      if(!TI && D) (posedge CP => (QN +: TE)) = (`F_FD1SHSP_CP_R_QN_R, `F_FD1SHSP_CP_R_QN_F);

	$setuphold(posedge CP &&& XorDTI_, posedge TE, `F_FD1SHSP_TE_CP_SETUP_posedge_posedge, `F_FD1SHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& XorDTI_, negedge TE, `F_FD1SHSP_TE_CP_SETUP_negedge_posedge, `F_FD1SHSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `F_FD1SHSP_TI_CP_SETUP_posedge_posedge, `F_FD1SHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `F_FD1SHSP_TI_CP_SETUP_negedge_posedge, `F_FD1SHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TEX, posedge D, `F_FD1SHSP_D_CP_SETUP_posedge_posedge, `F_FD1SHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TEX, negedge D, `F_FD1SHSP_D_CP_SETUP_negedge_posedge, `F_FD1SHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `F_FD1SHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `F_FD1SHSP_CP_PWH, 0, Notifier);
`else
     (posedge CP => (Q +: Mux21DTITE_)) = (`F_FD1SHSP_CP_R_Q_R, `F_FD1SHSP_CP_R_Q_F);
     (posedge CP => (QN -: Mux21DTITE_)) = (`F_FD1SHSP_CP_R_QN_R, `F_FD1SHSP_CP_R_QN_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `F_FD1SHSP_TE_CP_SETUP_posedge_posedge, `F_FD1SHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `F_FD1SHSP_TE_CP_SETUP_negedge_posedge, `F_FD1SHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `F_FD1SHSP_TI_CP_SETUP_posedge_posedge, `F_FD1SHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `F_FD1SHSP_TI_CP_SETUP_negedge_posedge, `F_FD1SHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `F_FD1SHSP_D_CP_SETUP_posedge_posedge, `F_FD1SHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `F_FD1SHSP_D_CP_SETUP_negedge_posedge, `F_FD1SHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `F_FD1SHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `F_FD1SHSP_CP_PWH, 0, Notifier);
`endif 
   endspecify
`endif


endmodule // F_FD1SHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:07 and Version :1.1 //
 
//  START 

// CELL FD1SQHS
 
`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 
 
`define FD1SQHS_CP_R_Q_R 0.1
`define FD1SQHS_CP_R_Q_F 0.1
`define FD1SQHS_CP_PWH 0.1
`define FD1SQHS_CP_PWL 0.1
`define FD1SQHS_D_CP_SETUP_posedge_posedge 0.1
`define FD1SQHS_D_CP_SETUP_negedge_posedge 0.1
`define FD1SQHS_D_CP_HOLD_posedge_posedge 0.1
`define FD1SQHS_D_CP_HOLD_negedge_posedge 0.1
`define FD1SQHS_TI_CP_SETUP_posedge_posedge 0.1
`define FD1SQHS_TI_CP_SETUP_negedge_posedge 0.1
`define FD1SQHS_TI_CP_HOLD_posedge_posedge 0.1
`define FD1SQHS_TI_CP_HOLD_negedge_posedge 0.1
`define FD1SQHS_TE_CP_SETUP_posedge_posedge 0.1
`define FD1SQHS_TE_CP_SETUP_negedge_posedge 0.1
`define FD1SQHS_TE_CP_HOLD_posedge_posedge 0.1
`define FD1SQHS_TE_CP_HOLD_negedge_posedge 0.1
 
module FD1SQHS (Q, D, CP, TI, TE);
 
   output Q;
   input D;
   input CP;
   input TI;
   input TE;
 
   reg Notifier;
 
   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);
 
   U_FD_P_NOTI u1 (IQ, Mux21DTITE_, CP, Notifier);
 
   buf  u2 (Q, IQ);
 
 
 
`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault
      if(!TE) (posedge CP => (Q +: D)) = (`FD1SQHS_CP_R_Q_R, `FD1SQHS_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD1SQHS_CP_R_Q_R, `FD1SQHS_CP_R_Q_F);
      if(!D && TI) (posedge CP => (Q +: TE)) = (`FD1SQHS_CP_R_Q_R, `FD1SQHS_CP_R_Q_F);
      if(!TI && D) (posedge CP => (Q -: TE)) = (`FD1SQHS_CP_R_Q_R, `FD1SQHS_CP_R_Q_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `FD1SQHS_TE_CP_SETUP_posedge_posedge, `FD1SQHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `FD1SQHS_TE_CP_SETUP_negedge_posedge, `FD1SQHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD1SQHS_TI_CP_SETUP_posedge_posedge, `FD1SQHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD1SQHS_TI_CP_SETUP_negedge_posedge, `FD1SQHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `FD1SQHS_D_CP_SETUP_posedge_posedge, `FD1SQHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `FD1SQHS_D_CP_SETUP_negedge_posedge, `FD1SQHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD1SQHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1SQHS_CP_PWH, 0, Notifier);
`else
     (posedge CP => (Q +: Mux21DTITE_)) = (`FD1SQHS_CP_R_Q_R, `FD1SQHS_CP_R_Q_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `FD1SQHS_TE_CP_SETUP_posedge_posedge, `FD1SQHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `FD1SQHS_TE_CP_SETUP_negedge_posedge, `FD1SQHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD1SQHS_TI_CP_SETUP_posedge_posedge, `FD1SQHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD1SQHS_TI_CP_SETUP_negedge_posedge, `FD1SQHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `FD1SQHS_D_CP_SETUP_posedge_posedge, `FD1SQHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `FD1SQHS_D_CP_SETUP_negedge_posedge, `FD1SQHS_D_CP_HOLD_negedge_posedge, Notifier);
      $width(negedge CP, `FD1SQHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1SQHS_CP_PWH, 0, Notifier);
`endif
   endspecify
`endif
 
 
endmodule // FD1SQHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
 
//  END
// Created from CVS on Date :1998/07/07 13:15:09 and Version :1.1 //
 
//  START
 





// CELL FD1SQHSP
 
`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 
 
`define FD1SQHSP_CP_R_Q_R 0.1
`define FD1SQHSP_CP_R_Q_F 0.1
`define FD1SQHSP_CP_PWH 0.1
`define FD1SQHSP_CP_PWL 0.1
`define FD1SQHSP_D_CP_SETUP_posedge_posedge 0.1
`define FD1SQHSP_D_CP_SETUP_negedge_posedge 0.1
`define FD1SQHSP_D_CP_HOLD_posedge_posedge 0.1
`define FD1SQHSP_D_CP_HOLD_negedge_posedge 0.1
`define FD1SQHSP_TI_CP_SETUP_posedge_posedge 0.1
`define FD1SQHSP_TI_CP_SETUP_negedge_posedge 0.1
`define FD1SQHSP_TI_CP_HOLD_posedge_posedge 0.1
`define FD1SQHSP_TI_CP_HOLD_negedge_posedge 0.1
`define FD1SQHSP_TE_CP_SETUP_posedge_posedge 0.1
`define FD1SQHSP_TE_CP_SETUP_negedge_posedge 0.1
`define FD1SQHSP_TE_CP_HOLD_posedge_posedge 0.1
`define FD1SQHSP_TE_CP_HOLD_negedge_posedge 0.1
 
module FD1SQHSP (Q, D, CP, TI, TE);
 
   output Q;
   input D;
   input CP;
   input TI;
   input TE;
 
   reg Notifier;
 
   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);
 
   U_FD_P_NOTI u1 (IQ, Mux21DTITE_, CP, Notifier);
 
   buf  u2 (Q, IQ);
 
 
 
`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault
      if(!TE) (posedge CP => (Q +: D)) = (`FD1SQHSP_CP_R_Q_R, `FD1SQHSP_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD1SQHSP_CP_R_Q_R, `FD1SQHSP_CP_R_Q_F);
      if(!D && TI) (posedge CP => (Q +: TE)) = (`FD1SQHSP_CP_R_Q_R, `FD1SQHSP_CP_R_Q_F);
      if(!TI && D) (posedge CP => (Q -: TE)) = (`FD1SQHSP_CP_R_Q_R, `FD1SQHSP_CP_R_Q_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `FD1SQHSP_TE_CP_SETUP_posedge_posedge, `FD1SQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `FD1SQHSP_TE_CP_SETUP_negedge_posedge, `FD1SQHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD1SQHSP_TI_CP_SETUP_posedge_posedge, `FD1SQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD1SQHSP_TI_CP_SETUP_negedge_posedge, `FD1SQHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `FD1SQHSP_D_CP_SETUP_posedge_posedge, `FD1SQHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `FD1SQHSP_D_CP_SETUP_negedge_posedge, `FD1SQHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD1SQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1SQHSP_CP_PWH, 0, Notifier);
`else
     (posedge CP => (Q +: Mux21DTITE_)) = (`FD1SQHSP_CP_R_Q_R, `FD1SQHSP_CP_R_Q_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `FD1SQHSP_TE_CP_SETUP_posedge_posedge, `FD1SQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `FD1SQHSP_TE_CP_SETUP_negedge_posedge, `FD1SQHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD1SQHSP_TI_CP_SETUP_posedge_posedge, `FD1SQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD1SQHSP_TI_CP_SETUP_negedge_posedge, `FD1SQHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `FD1SQHSP_D_CP_SETUP_posedge_posedge, `FD1SQHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `FD1SQHSP_D_CP_SETUP_negedge_posedge, `FD1SQHSP_D_CP_HOLD_negedge_posedge, Notifier);
      $width(negedge CP, `FD1SQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1SQHSP_CP_PWH, 0, Notifier);
`endif
   endspecify
`endif
 
 
endmodule // FD1SQHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
 
//  END
// Created from CVS on Date :1998/07/07 13:15:09 and Version :1.1 //
 
//  START
 





// CELL FD1SQHSX4
 
`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 
 
`define FD1SQHSX4_CP_R_Q_R 0.1
`define FD1SQHSX4_CP_R_Q_F 0.1
`define FD1SQHSX4_CP_PWH 0.1
`define FD1SQHSX4_CP_PWL 0.1
`define FD1SQHSX4_D_CP_SETUP_posedge_posedge 0.1
`define FD1SQHSX4_D_CP_SETUP_negedge_posedge 0.1
`define FD1SQHSX4_D_CP_HOLD_posedge_posedge 0.1
`define FD1SQHSX4_D_CP_HOLD_negedge_posedge 0.1
`define FD1SQHSX4_TI_CP_SETUP_posedge_posedge 0.1
`define FD1SQHSX4_TI_CP_SETUP_negedge_posedge 0.1
`define FD1SQHSX4_TI_CP_HOLD_posedge_posedge 0.1
`define FD1SQHSX4_TI_CP_HOLD_negedge_posedge 0.1
`define FD1SQHSX4_TE_CP_SETUP_posedge_posedge 0.1
`define FD1SQHSX4_TE_CP_SETUP_negedge_posedge 0.1
`define FD1SQHSX4_TE_CP_HOLD_posedge_posedge 0.1
`define FD1SQHSX4_TE_CP_HOLD_negedge_posedge 0.1
 
module FD1SQHSX4 (Q, D, CP, TI, TE);
 
   output Q;
   input D;
   input CP;
   input TI;
   input TE;
 
   reg Notifier;
 
   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);
 
   U_FD_P_NOTI u1 (IQ, Mux21DTITE_, CP, Notifier);
 
   buf  u2 (Q, IQ);
 
 
 
`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault
      if(!TE) (posedge CP => (Q +: D)) = (`FD1SQHSX4_CP_R_Q_R, `FD1SQHSX4_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD1SQHSX4_CP_R_Q_R, `FD1SQHSX4_CP_R_Q_F);
      if(!D && TI) (posedge CP => (Q +: TE)) = (`FD1SQHSX4_CP_R_Q_R, `FD1SQHSX4_CP_R_Q_F);
      if(!TI && D) (posedge CP => (Q -: TE)) = (`FD1SQHSX4_CP_R_Q_R, `FD1SQHSX4_CP_R_Q_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `FD1SQHSX4_TE_CP_SETUP_posedge_posedge, `FD1SQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `FD1SQHSX4_TE_CP_SETUP_negedge_posedge, `FD1SQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD1SQHSX4_TI_CP_SETUP_posedge_posedge, `FD1SQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD1SQHSX4_TI_CP_SETUP_negedge_posedge, `FD1SQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `FD1SQHSX4_D_CP_SETUP_posedge_posedge, `FD1SQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `FD1SQHSX4_D_CP_SETUP_negedge_posedge, `FD1SQHSX4_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD1SQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1SQHSX4_CP_PWH, 0, Notifier);
`else
     (posedge CP => (Q +: Mux21DTITE_)) = (`FD1SQHSX4_CP_R_Q_R, `FD1SQHSX4_CP_R_Q_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `FD1SQHSX4_TE_CP_SETUP_posedge_posedge, `FD1SQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `FD1SQHSX4_TE_CP_SETUP_negedge_posedge, `FD1SQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD1SQHSX4_TI_CP_SETUP_posedge_posedge, `FD1SQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD1SQHSX4_TI_CP_SETUP_negedge_posedge, `FD1SQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `FD1SQHSX4_D_CP_SETUP_posedge_posedge, `FD1SQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `FD1SQHSX4_D_CP_SETUP_negedge_posedge, `FD1SQHSX4_D_CP_HOLD_negedge_posedge, Notifier);
      $width(negedge CP, `FD1SQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1SQHSX4_CP_PWH, 0, Notifier);
`endif
   endspecify
`endif
 
 
endmodule // FD1SQHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
 
//  END
// Created from CVS on Date :1998/07/07 13:15:09 and Version :1.1 //
 
//  START
 





// CELL FDM1SQHS
 
`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 
 
`define FDM1SQHS_CP_R_Q_R 0.1
`define FDM1SQHS_CP_R_Q_F 0.1
`define FDM1SQHS_CP_PWH 0.1
`define FDM1SQHS_CP_PWL 0.1
`define FDM1SQHS_D_CP_SETUP_posedge_posedge 0.1
`define FDM1SQHS_D_CP_SETUP_negedge_posedge 0.1
`define FDM1SQHS_D_CP_HOLD_posedge_posedge 0.1
`define FDM1SQHS_D_CP_HOLD_negedge_posedge 0.1
`define FDM1SQHS_TI_CP_SETUP_posedge_posedge 0.1
`define FDM1SQHS_TI_CP_SETUP_negedge_posedge 0.1
`define FDM1SQHS_TI_CP_HOLD_posedge_posedge 0.1
`define FDM1SQHS_TI_CP_HOLD_negedge_posedge 0.1
`define FDM1SQHS_TE_CP_SETUP_posedge_posedge 0.1
`define FDM1SQHS_TE_CP_SETUP_negedge_posedge 0.1
`define FDM1SQHS_TE_CP_HOLD_posedge_posedge 0.1
`define FDM1SQHS_TE_CP_HOLD_negedge_posedge 0.1
 
module FDM1SQHS (Q, D, CP, TI, TE);
 
   output Q;
   input D;
   input CP;
   input TI;
   input TE;
 
   reg Notifier;
 
   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);
 
   U_FD_P_NOTI u1 (IQ, Mux21DTITE_, CP, Notifier);
 
   buf  u2 (Q, IQ);
 
 
 
`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault
      if(!TE) (posedge CP => (Q +: D)) = (`FDM1SQHS_CP_R_Q_R, `FDM1SQHS_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FDM1SQHS_CP_R_Q_R, `FDM1SQHS_CP_R_Q_F);
      if(!D && TI) (posedge CP => (Q +: TE)) = (`FDM1SQHS_CP_R_Q_R, `FDM1SQHS_CP_R_Q_F);
      if(!TI && D) (posedge CP => (Q -: TE)) = (`FDM1SQHS_CP_R_Q_R, `FDM1SQHS_CP_R_Q_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `FDM1SQHS_TE_CP_SETUP_posedge_posedge, `FDM1SQHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `FDM1SQHS_TE_CP_SETUP_negedge_posedge, `FDM1SQHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FDM1SQHS_TI_CP_SETUP_posedge_posedge, `FDM1SQHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FDM1SQHS_TI_CP_SETUP_negedge_posedge, `FDM1SQHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `FDM1SQHS_D_CP_SETUP_posedge_posedge, `FDM1SQHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `FDM1SQHS_D_CP_SETUP_negedge_posedge, `FDM1SQHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDM1SQHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FDM1SQHS_CP_PWH, 0, Notifier);
`else
     (posedge CP => (Q +: Mux21DTITE_)) = (`FDM1SQHS_CP_R_Q_R, `FDM1SQHS_CP_R_Q_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `FDM1SQHS_TE_CP_SETUP_posedge_posedge, `FDM1SQHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `FDM1SQHS_TE_CP_SETUP_negedge_posedge, `FDM1SQHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FDM1SQHS_TI_CP_SETUP_posedge_posedge, `FDM1SQHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FDM1SQHS_TI_CP_SETUP_negedge_posedge, `FDM1SQHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `FDM1SQHS_D_CP_SETUP_posedge_posedge, `FDM1SQHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `FDM1SQHS_D_CP_SETUP_negedge_posedge, `FDM1SQHS_D_CP_HOLD_negedge_posedge, Notifier);
      $width(negedge CP, `FDM1SQHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FDM1SQHS_CP_PWH, 0, Notifier);
`endif
   endspecify
`endif
 
 
endmodule // FDM1SQHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
 
//  END
// Created from CVS on Date :1998/07/07 13:15:09 and Version :1.1 //
 
//  START
 





// CELL FDM1SQHSP
 
`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 
 
`define FDM1SQHSP_CP_R_Q_R 0.1
`define FDM1SQHSP_CP_R_Q_F 0.1
`define FDM1SQHSP_CP_PWH 0.1
`define FDM1SQHSP_CP_PWL 0.1
`define FDM1SQHSP_D_CP_SETUP_posedge_posedge 0.1
`define FDM1SQHSP_D_CP_SETUP_negedge_posedge 0.1
`define FDM1SQHSP_D_CP_HOLD_posedge_posedge 0.1
`define FDM1SQHSP_D_CP_HOLD_negedge_posedge 0.1
`define FDM1SQHSP_TI_CP_SETUP_posedge_posedge 0.1
`define FDM1SQHSP_TI_CP_SETUP_negedge_posedge 0.1
`define FDM1SQHSP_TI_CP_HOLD_posedge_posedge 0.1
`define FDM1SQHSP_TI_CP_HOLD_negedge_posedge 0.1
`define FDM1SQHSP_TE_CP_SETUP_posedge_posedge 0.1
`define FDM1SQHSP_TE_CP_SETUP_negedge_posedge 0.1
`define FDM1SQHSP_TE_CP_HOLD_posedge_posedge 0.1
`define FDM1SQHSP_TE_CP_HOLD_negedge_posedge 0.1
 
module FDM1SQHSP (Q, D, CP, TI, TE);
 
   output Q;
   input D;
   input CP;
   input TI;
   input TE;
 
   reg Notifier;
 
   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);
 
   U_FD_P_NOTI u1 (IQ, Mux21DTITE_, CP, Notifier);
 
   buf  u2 (Q, IQ);
 
 
 
`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault
      if(!TE) (posedge CP => (Q +: D)) = (`FDM1SQHSP_CP_R_Q_R, `FDM1SQHSP_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FDM1SQHSP_CP_R_Q_R, `FDM1SQHSP_CP_R_Q_F);
      if(!D && TI) (posedge CP => (Q +: TE)) = (`FDM1SQHSP_CP_R_Q_R, `FDM1SQHSP_CP_R_Q_F);
      if(!TI && D) (posedge CP => (Q -: TE)) = (`FDM1SQHSP_CP_R_Q_R, `FDM1SQHSP_CP_R_Q_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `FDM1SQHSP_TE_CP_SETUP_posedge_posedge, `FDM1SQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `FDM1SQHSP_TE_CP_SETUP_negedge_posedge, `FDM1SQHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FDM1SQHSP_TI_CP_SETUP_posedge_posedge, `FDM1SQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FDM1SQHSP_TI_CP_SETUP_negedge_posedge, `FDM1SQHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `FDM1SQHSP_D_CP_SETUP_posedge_posedge, `FDM1SQHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `FDM1SQHSP_D_CP_SETUP_negedge_posedge, `FDM1SQHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDM1SQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FDM1SQHSP_CP_PWH, 0, Notifier);
`else
     (posedge CP => (Q +: Mux21DTITE_)) = (`FDM1SQHSP_CP_R_Q_R, `FDM1SQHSP_CP_R_Q_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `FDM1SQHSP_TE_CP_SETUP_posedge_posedge, `FDM1SQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `FDM1SQHSP_TE_CP_SETUP_negedge_posedge, `FDM1SQHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FDM1SQHSP_TI_CP_SETUP_posedge_posedge, `FDM1SQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FDM1SQHSP_TI_CP_SETUP_negedge_posedge, `FDM1SQHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `FDM1SQHSP_D_CP_SETUP_posedge_posedge, `FDM1SQHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `FDM1SQHSP_D_CP_SETUP_negedge_posedge, `FDM1SQHSP_D_CP_HOLD_negedge_posedge, Notifier);
      $width(negedge CP, `FDM1SQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FDM1SQHSP_CP_PWH, 0, Notifier);
`endif
   endspecify
`endif
 
 
endmodule // FDM1SQHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
 
//  END
// Created from CVS on Date :1998/07/07 13:15:09 and Version :1.1 //
 
//  START
 





// CELL F_FD1SQHS
 
`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 
 
`define F_FD1SQHS_CP_R_Q_R 0.1
`define F_FD1SQHS_CP_R_Q_F 0.1
`define F_FD1SQHS_CP_PWH 0.1
`define F_FD1SQHS_CP_PWL 0.1
`define F_FD1SQHS_D_CP_SETUP_posedge_posedge 0.1
`define F_FD1SQHS_D_CP_SETUP_negedge_posedge 0.1
`define F_FD1SQHS_D_CP_HOLD_posedge_posedge 0.1
`define F_FD1SQHS_D_CP_HOLD_negedge_posedge 0.1
`define F_FD1SQHS_TI_CP_SETUP_posedge_posedge 0.1
`define F_FD1SQHS_TI_CP_SETUP_negedge_posedge 0.1
`define F_FD1SQHS_TI_CP_HOLD_posedge_posedge 0.1
`define F_FD1SQHS_TI_CP_HOLD_negedge_posedge 0.1
`define F_FD1SQHS_TE_CP_SETUP_posedge_posedge 0.1
`define F_FD1SQHS_TE_CP_SETUP_negedge_posedge 0.1
`define F_FD1SQHS_TE_CP_HOLD_posedge_posedge 0.1
`define F_FD1SQHS_TE_CP_HOLD_negedge_posedge 0.1
 
module F_FD1SQHS (Q, D, CP, TI, TE);
 
   output Q;
   input D;
   input CP;
   input TI;
   input TE;
 
   reg Notifier;
 
   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);
 
   U_FD_P_NOTI u1 (IQ, Mux21DTITE_, CP, Notifier);
 
   buf  u2 (Q, IQ);
 
 
 
`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault
      if(!TE) (posedge CP => (Q +: D)) = (`F_FD1SQHS_CP_R_Q_R, `F_FD1SQHS_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`F_FD1SQHS_CP_R_Q_R, `F_FD1SQHS_CP_R_Q_F);
      if(!D && TI) (posedge CP => (Q +: TE)) = (`F_FD1SQHS_CP_R_Q_R, `F_FD1SQHS_CP_R_Q_F);
      if(!TI && D) (posedge CP => (Q -: TE)) = (`F_FD1SQHS_CP_R_Q_R, `F_FD1SQHS_CP_R_Q_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `F_FD1SQHS_TE_CP_SETUP_posedge_posedge, `F_FD1SQHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `F_FD1SQHS_TE_CP_SETUP_negedge_posedge, `F_FD1SQHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `F_FD1SQHS_TI_CP_SETUP_posedge_posedge, `F_FD1SQHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `F_FD1SQHS_TI_CP_SETUP_negedge_posedge, `F_FD1SQHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `F_FD1SQHS_D_CP_SETUP_posedge_posedge, `F_FD1SQHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `F_FD1SQHS_D_CP_SETUP_negedge_posedge, `F_FD1SQHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `F_FD1SQHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `F_FD1SQHS_CP_PWH, 0, Notifier);
`else
     (posedge CP => (Q +: Mux21DTITE_)) = (`F_FD1SQHS_CP_R_Q_R, `F_FD1SQHS_CP_R_Q_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `F_FD1SQHS_TE_CP_SETUP_posedge_posedge, `F_FD1SQHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `F_FD1SQHS_TE_CP_SETUP_negedge_posedge, `F_FD1SQHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `F_FD1SQHS_TI_CP_SETUP_posedge_posedge, `F_FD1SQHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `F_FD1SQHS_TI_CP_SETUP_negedge_posedge, `F_FD1SQHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `F_FD1SQHS_D_CP_SETUP_posedge_posedge, `F_FD1SQHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `F_FD1SQHS_D_CP_SETUP_negedge_posedge, `F_FD1SQHS_D_CP_HOLD_negedge_posedge, Notifier);
      $width(negedge CP, `F_FD1SQHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `F_FD1SQHS_CP_PWH, 0, Notifier);
`endif
   endspecify
`endif
 
 
endmodule // F_FD1SQHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
 
//  END
// Created from CVS on Date :1998/07/07 13:15:09 and Version :1.1 //
 
//  START
 





// CELL F_FD1SQHSP
 
`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 
 
`define F_FD1SQHSP_CP_R_Q_R 0.1
`define F_FD1SQHSP_CP_R_Q_F 0.1
`define F_FD1SQHSP_CP_PWH 0.1
`define F_FD1SQHSP_CP_PWL 0.1
`define F_FD1SQHSP_D_CP_SETUP_posedge_posedge 0.1
`define F_FD1SQHSP_D_CP_SETUP_negedge_posedge 0.1
`define F_FD1SQHSP_D_CP_HOLD_posedge_posedge 0.1
`define F_FD1SQHSP_D_CP_HOLD_negedge_posedge 0.1
`define F_FD1SQHSP_TI_CP_SETUP_posedge_posedge 0.1
`define F_FD1SQHSP_TI_CP_SETUP_negedge_posedge 0.1
`define F_FD1SQHSP_TI_CP_HOLD_posedge_posedge 0.1
`define F_FD1SQHSP_TI_CP_HOLD_negedge_posedge 0.1
`define F_FD1SQHSP_TE_CP_SETUP_posedge_posedge 0.1
`define F_FD1SQHSP_TE_CP_SETUP_negedge_posedge 0.1
`define F_FD1SQHSP_TE_CP_HOLD_posedge_posedge 0.1
`define F_FD1SQHSP_TE_CP_HOLD_negedge_posedge 0.1
 
module F_FD1SQHSP (Q, D, CP, TI, TE);
 
   output Q;
   input D;
   input CP;
   input TI;
   input TE;
 
   reg Notifier;
 
   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);
 
   U_FD_P_NOTI u1 (IQ, Mux21DTITE_, CP, Notifier);
 
   buf  u2 (Q, IQ);
 
 
 
`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault
      if(!TE) (posedge CP => (Q +: D)) = (`F_FD1SQHSP_CP_R_Q_R, `F_FD1SQHSP_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`F_FD1SQHSP_CP_R_Q_R, `F_FD1SQHSP_CP_R_Q_F);
      if(!D && TI) (posedge CP => (Q +: TE)) = (`F_FD1SQHSP_CP_R_Q_R, `F_FD1SQHSP_CP_R_Q_F);
      if(!TI && D) (posedge CP => (Q -: TE)) = (`F_FD1SQHSP_CP_R_Q_R, `F_FD1SQHSP_CP_R_Q_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `F_FD1SQHSP_TE_CP_SETUP_posedge_posedge, `F_FD1SQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `F_FD1SQHSP_TE_CP_SETUP_negedge_posedge, `F_FD1SQHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `F_FD1SQHSP_TI_CP_SETUP_posedge_posedge, `F_FD1SQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `F_FD1SQHSP_TI_CP_SETUP_negedge_posedge, `F_FD1SQHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `F_FD1SQHSP_D_CP_SETUP_posedge_posedge, `F_FD1SQHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `F_FD1SQHSP_D_CP_SETUP_negedge_posedge, `F_FD1SQHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `F_FD1SQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `F_FD1SQHSP_CP_PWH, 0, Notifier);
`else
     (posedge CP => (Q +: Mux21DTITE_)) = (`F_FD1SQHSP_CP_R_Q_R, `F_FD1SQHSP_CP_R_Q_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `F_FD1SQHSP_TE_CP_SETUP_posedge_posedge, `F_FD1SQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `F_FD1SQHSP_TE_CP_SETUP_negedge_posedge, `F_FD1SQHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `F_FD1SQHSP_TI_CP_SETUP_posedge_posedge, `F_FD1SQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `F_FD1SQHSP_TI_CP_SETUP_negedge_posedge, `F_FD1SQHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `F_FD1SQHSP_D_CP_SETUP_posedge_posedge, `F_FD1SQHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `F_FD1SQHSP_D_CP_SETUP_negedge_posedge, `F_FD1SQHSP_D_CP_HOLD_negedge_posedge, Notifier);
      $width(negedge CP, `F_FD1SQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `F_FD1SQHSP_CP_PWH, 0, Notifier);
`endif
   endspecify
`endif
 
 
endmodule // F_FD1SQHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
 
//  END
// Created from CVS on Date :1998/07/07 13:15:09 and Version :1.1 //
 
//  START
 





// CELL F_FD1SQHSX4
 
`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 
 
`define F_FD1SQHSX4_CP_R_Q_R 0.1
`define F_FD1SQHSX4_CP_R_Q_F 0.1
`define F_FD1SQHSX4_CP_PWH 0.1
`define F_FD1SQHSX4_CP_PWL 0.1
`define F_FD1SQHSX4_D_CP_SETUP_posedge_posedge 0.1
`define F_FD1SQHSX4_D_CP_SETUP_negedge_posedge 0.1
`define F_FD1SQHSX4_D_CP_HOLD_posedge_posedge 0.1
`define F_FD1SQHSX4_D_CP_HOLD_negedge_posedge 0.1
`define F_FD1SQHSX4_TI_CP_SETUP_posedge_posedge 0.1
`define F_FD1SQHSX4_TI_CP_SETUP_negedge_posedge 0.1
`define F_FD1SQHSX4_TI_CP_HOLD_posedge_posedge 0.1
`define F_FD1SQHSX4_TI_CP_HOLD_negedge_posedge 0.1
`define F_FD1SQHSX4_TE_CP_SETUP_posedge_posedge 0.1
`define F_FD1SQHSX4_TE_CP_SETUP_negedge_posedge 0.1
`define F_FD1SQHSX4_TE_CP_HOLD_posedge_posedge 0.1
`define F_FD1SQHSX4_TE_CP_HOLD_negedge_posedge 0.1
 
module F_FD1SQHSX4 (Q, D, CP, TI, TE);
 
   output Q;
   input D;
   input CP;
   input TI;
   input TE;
 
   reg Notifier;
 
   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);
 
   U_FD_P_NOTI u1 (IQ, Mux21DTITE_, CP, Notifier);
 
   buf  u2 (Q, IQ);
 
 
 
`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault
      if(!TE) (posedge CP => (Q +: D)) = (`F_FD1SQHSX4_CP_R_Q_R, `F_FD1SQHSX4_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`F_FD1SQHSX4_CP_R_Q_R, `F_FD1SQHSX4_CP_R_Q_F);
      if(!D && TI) (posedge CP => (Q +: TE)) = (`F_FD1SQHSX4_CP_R_Q_R, `F_FD1SQHSX4_CP_R_Q_F);
      if(!TI && D) (posedge CP => (Q -: TE)) = (`F_FD1SQHSX4_CP_R_Q_R, `F_FD1SQHSX4_CP_R_Q_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `F_FD1SQHSX4_TE_CP_SETUP_posedge_posedge, `F_FD1SQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `F_FD1SQHSX4_TE_CP_SETUP_negedge_posedge, `F_FD1SQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `F_FD1SQHSX4_TI_CP_SETUP_posedge_posedge, `F_FD1SQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `F_FD1SQHSX4_TI_CP_SETUP_negedge_posedge, `F_FD1SQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `F_FD1SQHSX4_D_CP_SETUP_posedge_posedge, `F_FD1SQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `F_FD1SQHSX4_D_CP_SETUP_negedge_posedge, `F_FD1SQHSX4_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `F_FD1SQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP, `F_FD1SQHSX4_CP_PWH, 0, Notifier);
`else
     (posedge CP => (Q +: Mux21DTITE_)) = (`F_FD1SQHSX4_CP_R_Q_R, `F_FD1SQHSX4_CP_R_Q_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `F_FD1SQHSX4_TE_CP_SETUP_posedge_posedge, `F_FD1SQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `F_FD1SQHSX4_TE_CP_SETUP_negedge_posedge, `F_FD1SQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `F_FD1SQHSX4_TI_CP_SETUP_posedge_posedge, `F_FD1SQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `F_FD1SQHSX4_TI_CP_SETUP_negedge_posedge, `F_FD1SQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `F_FD1SQHSX4_D_CP_SETUP_posedge_posedge, `F_FD1SQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `F_FD1SQHSX4_D_CP_SETUP_negedge_posedge, `F_FD1SQHSX4_D_CP_HOLD_negedge_posedge, Notifier);
      $width(negedge CP, `F_FD1SQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP, `F_FD1SQHSX4_CP_PWH, 0, Notifier);
`endif
   endspecify
`endif
 
 
endmodule // F_FD1SQHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
 
//  END
// Created from CVS on Date :1998/07/07 13:15:09 and Version :1.1 //
 
//  START
 





// CELL FD1THS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD1THS_CP_R_SO_R 0.1
`define FD1THS_CP_R_SO_F 0.1
`define FD1THS_CP_R_QN_F 0.1
`define FD1THS_CP_R_QN_R 0.1
`define FD1THS_CP_R_Q_R 0.1
`define FD1THS_CP_R_Q_F 0.1
`define FD1THS_CP_PWH 0.1
`define FD1THS_CP_PWL 0.1
`define FD1THS_D_CP_SETUP_posedge_posedge 0.1
`define FD1THS_D_CP_SETUP_negedge_posedge 0.1
`define FD1THS_D_CP_HOLD_posedge_posedge 0.1
`define FD1THS_D_CP_HOLD_negedge_posedge 0.1
`define FD1THS_TI_CP_SETUP_posedge_posedge 0.1
`define FD1THS_TI_CP_SETUP_negedge_posedge 0.1
`define FD1THS_TI_CP_HOLD_posedge_posedge 0.1
`define FD1THS_TI_CP_HOLD_negedge_posedge 0.1
`define FD1THS_TE_CP_SETUP_posedge_posedge 0.1
`define FD1THS_TE_CP_SETUP_negedge_posedge 0.1
`define FD1THS_TE_CP_HOLD_posedge_posedge 0.1
`define FD1THS_TE_CP_HOLD_negedge_posedge 0.1

module FD1THS (Q, QN, SO, D, CP, TI, TE);

   output Q;
   output QN;
   output SO;
   input D;
   input CP;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, Notifier);

   buf  u2 (Q, IQ);
   buf  u3 (SO, IQ);
   not  u4 (QN, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault

      if(!TE) (posedge CP => (Q +: D)) = (`FD1THS_CP_R_Q_R, `FD1THS_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD1THS_CP_R_Q_R, `FD1THS_CP_R_Q_F);
      if(!D && TI) (posedge CP => (Q +: TE)) = (`FD1THS_CP_R_Q_R, `FD1THS_CP_R_Q_F);
      if(!TI && D) (posedge CP => (Q -: TE)) = (`FD1THS_CP_R_Q_R, `FD1THS_CP_R_Q_F);
      if(!TE) (posedge CP => (QN -: D)) = (`FD1THS_CP_R_QN_R, `FD1THS_CP_R_QN_F);
      if(TE) (posedge CP => (QN -: TI)) = (`FD1THS_CP_R_QN_R, `FD1THS_CP_R_QN_F);
      if(!D && TI) (posedge CP => (QN -: TE)) = (`FD1THS_CP_R_QN_R, `FD1THS_CP_R_QN_F);
      if(!TI && D) (posedge CP => (QN +: TE)) = (`FD1THS_CP_R_QN_R, `FD1THS_CP_R_QN_F);
      if(!TE) (posedge CP => (SO +: D)) = (`FD1THS_CP_R_SO_R, `FD1THS_CP_R_SO_F);
      if(TE) (posedge CP => (SO +: TI)) = (`FD1THS_CP_R_SO_R, `FD1THS_CP_R_SO_F);
      if(!D && TI) (posedge CP => (SO +: TE)) = (`FD1THS_CP_R_SO_R, `FD1THS_CP_R_SO_F);
      if(!TI && D) (posedge CP => (SO -: TE)) = (`FD1THS_CP_R_SO_R, `FD1THS_CP_R_SO_F);

	$setuphold(posedge CP &&& XorDTI_, posedge TE, `FD1THS_TE_CP_SETUP_posedge_posedge, `FD1THS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& XorDTI_, negedge TE, `FD1THS_TE_CP_SETUP_negedge_posedge, `FD1THS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FD1THS_TI_CP_SETUP_posedge_posedge, `FD1THS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FD1THS_TI_CP_SETUP_negedge_posedge, `FD1THS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TEX, posedge D, `FD1THS_D_CP_SETUP_posedge_posedge, `FD1THS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TEX, negedge D, `FD1THS_D_CP_SETUP_negedge_posedge, `FD1THS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD1THS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1THS_CP_PWH, 0, Notifier);
`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FD1THS_CP_R_Q_R, `FD1THS_CP_R_Q_F);
      (posedge CP => (QN -: Mux21DTITE_)) = (`FD1THS_CP_R_QN_R, `FD1THS_CP_R_QN_F);
      (posedge CP => (SO +: Mux21DTITE_)) = (`FD1THS_CP_R_SO_R, `FD1THS_CP_R_SO_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `FD1THS_TE_CP_SETUP_posedge_posedge, `FD1THS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `FD1THS_TE_CP_SETUP_negedge_posedge, `FD1THS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD1THS_TI_CP_SETUP_posedge_posedge, `FD1THS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD1THS_TI_CP_SETUP_negedge_posedge, `FD1THS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `FD1THS_D_CP_SETUP_posedge_posedge, `FD1THS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `FD1THS_D_CP_SETUP_negedge_posedge, `FD1THS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD1THS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1THS_CP_PWH, 0, Notifier);

`endif
   endspecify
`endif


endmodule // FD1THS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:13 and Version :1.1 //
 
//  START 
// CELL FD1THSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD1THSP_CP_R_SO_R 0.1
`define FD1THSP_CP_R_SO_F 0.1
`define FD1THSP_CP_R_QN_F 0.1
`define FD1THSP_CP_R_QN_R 0.1
`define FD1THSP_CP_R_Q_R 0.1
`define FD1THSP_CP_R_Q_F 0.1
`define FD1THSP_CP_PWH 0.1
`define FD1THSP_CP_PWL 0.1
`define FD1THSP_D_CP_SETUP_posedge_posedge 0.1
`define FD1THSP_D_CP_SETUP_negedge_posedge 0.1
`define FD1THSP_D_CP_HOLD_posedge_posedge 0.1
`define FD1THSP_D_CP_HOLD_negedge_posedge 0.1
`define FD1THSP_TI_CP_SETUP_posedge_posedge 0.1
`define FD1THSP_TI_CP_SETUP_negedge_posedge 0.1
`define FD1THSP_TI_CP_HOLD_posedge_posedge 0.1
`define FD1THSP_TI_CP_HOLD_negedge_posedge 0.1
`define FD1THSP_TE_CP_SETUP_posedge_posedge 0.1
`define FD1THSP_TE_CP_SETUP_negedge_posedge 0.1
`define FD1THSP_TE_CP_HOLD_posedge_posedge 0.1
`define FD1THSP_TE_CP_HOLD_negedge_posedge 0.1

module FD1THSP (Q, QN, SO, D, CP, TI, TE);

   output Q;
   output QN;
   output SO;
   input D;
   input CP;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, Notifier);

   buf  u2 (Q, IQ);
   buf  u3 (SO, IQ);
   not  u4 (QN, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault

      if(!TE) (posedge CP => (Q +: D)) = (`FD1THSP_CP_R_Q_R, `FD1THSP_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD1THSP_CP_R_Q_R, `FD1THSP_CP_R_Q_F);
      if(!D && TI) (posedge CP => (Q +: TE)) = (`FD1THSP_CP_R_Q_R, `FD1THSP_CP_R_Q_F);
      if(!TI && D) (posedge CP => (Q -: TE)) = (`FD1THSP_CP_R_Q_R, `FD1THSP_CP_R_Q_F);
      if(!TE) (posedge CP => (QN -: D)) = (`FD1THSP_CP_R_QN_R, `FD1THSP_CP_R_QN_F);
      if(TE) (posedge CP => (QN -: TI)) = (`FD1THSP_CP_R_QN_R, `FD1THSP_CP_R_QN_F);
      if(!D && TI) (posedge CP => (QN -: TE)) = (`FD1THSP_CP_R_QN_R, `FD1THSP_CP_R_QN_F);
      if(!TI && D) (posedge CP => (QN +: TE)) = (`FD1THSP_CP_R_QN_R, `FD1THSP_CP_R_QN_F);
      if(!TE) (posedge CP => (SO +: D)) = (`FD1THSP_CP_R_SO_R, `FD1THSP_CP_R_SO_F);
      if(TE) (posedge CP => (SO +: TI)) = (`FD1THSP_CP_R_SO_R, `FD1THSP_CP_R_SO_F);
      if(!D && TI) (posedge CP => (SO +: TE)) = (`FD1THSP_CP_R_SO_R, `FD1THSP_CP_R_SO_F);
      if(!TI && D) (posedge CP => (SO -: TE)) = (`FD1THSP_CP_R_SO_R, `FD1THSP_CP_R_SO_F);

	$setuphold(posedge CP &&& XorDTI_, posedge TE, `FD1THSP_TE_CP_SETUP_posedge_posedge, `FD1THSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& XorDTI_, negedge TE, `FD1THSP_TE_CP_SETUP_negedge_posedge, `FD1THSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FD1THSP_TI_CP_SETUP_posedge_posedge, `FD1THSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FD1THSP_TI_CP_SETUP_negedge_posedge, `FD1THSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TEX, posedge D, `FD1THSP_D_CP_SETUP_posedge_posedge, `FD1THSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TEX, negedge D, `FD1THSP_D_CP_SETUP_negedge_posedge, `FD1THSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD1THSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1THSP_CP_PWH, 0, Notifier);
`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FD1THSP_CP_R_Q_R, `FD1THSP_CP_R_Q_F);
      (posedge CP => (QN -: Mux21DTITE_)) = (`FD1THSP_CP_R_QN_R, `FD1THSP_CP_R_QN_F);
      (posedge CP => (SO +: Mux21DTITE_)) = (`FD1THSP_CP_R_SO_R, `FD1THSP_CP_R_SO_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `FD1THSP_TE_CP_SETUP_posedge_posedge, `FD1THSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `FD1THSP_TE_CP_SETUP_negedge_posedge, `FD1THSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD1THSP_TI_CP_SETUP_posedge_posedge, `FD1THSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD1THSP_TI_CP_SETUP_negedge_posedge, `FD1THSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `FD1THSP_D_CP_SETUP_posedge_posedge, `FD1THSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `FD1THSP_D_CP_SETUP_negedge_posedge, `FD1THSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD1THSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1THSP_CP_PWH, 0, Notifier);

`endif
   endspecify
`endif


endmodule // FD1THSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:13 and Version :1.1 //
 
//  START 
// CELL FD1TQHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD1TQHS_CP_R_SO_R 0.1
`define FD1TQHS_CP_R_SO_F 0.1
`define FD1TQHS_CP_R_Q_R 0.1
`define FD1TQHS_CP_R_Q_F 0.1
`define FD1TQHS_CP_PWH 0.1
`define FD1TQHS_CP_PWL 0.1
`define FD1TQHS_D_CP_SETUP_posedge_posedge 0.1
`define FD1TQHS_D_CP_SETUP_negedge_posedge 0.1
`define FD1TQHS_D_CP_HOLD_posedge_posedge 0.1
`define FD1TQHS_D_CP_HOLD_negedge_posedge 0.1
`define FD1TQHS_TI_CP_SETUP_posedge_posedge 0.1
`define FD1TQHS_TI_CP_SETUP_negedge_posedge 0.1
`define FD1TQHS_TI_CP_HOLD_posedge_posedge 0.1
`define FD1TQHS_TI_CP_HOLD_negedge_posedge 0.1
`define FD1TQHS_TE_CP_SETUP_posedge_posedge 0.1
`define FD1TQHS_TE_CP_SETUP_negedge_posedge 0.1
`define FD1TQHS_TE_CP_HOLD_posedge_posedge 0.1
`define FD1TQHS_TE_CP_HOLD_negedge_posedge 0.1

module FD1TQHS (Q, SO, D, CP, TI, TE);

   output Q;
   output SO;
   input D;
   input CP;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, Notifier);

   buf  u2 (Q, IQ);
buf  u3 (SO, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault

      if(!TE) (posedge CP => (Q +: D)) = (`FD1TQHS_CP_R_Q_R, `FD1TQHS_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD1TQHS_CP_R_Q_R, `FD1TQHS_CP_R_Q_F);
      if(!D && TI) (posedge CP => (Q +: TE)) = (`FD1TQHS_CP_R_Q_R, `FD1TQHS_CP_R_Q_F);
      if(!TI && D) (posedge CP => (Q -: TE)) = (`FD1TQHS_CP_R_Q_R, `FD1TQHS_CP_R_Q_F);
      if(!TE) (posedge CP => (SO +: D)) = (`FD1TQHS_CP_R_SO_R, `FD1TQHS_CP_R_SO_F);
      if(TE) (posedge CP => (SO +: TI)) = (`FD1TQHS_CP_R_SO_R, `FD1TQHS_CP_R_SO_F);
      if(!D && TI) (posedge CP => (SO +: TE)) = (`FD1TQHS_CP_R_SO_R, `FD1TQHS_CP_R_SO_F);
      if(!TI && D) (posedge CP => (SO -: TE)) = (`FD1TQHS_CP_R_SO_R, `FD1TQHS_CP_R_SO_F);

	$setuphold(posedge CP &&& XorDTI_, posedge TE, `FD1TQHS_TE_CP_SETUP_posedge_posedge, `FD1TQHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& XorDTI_, negedge TE, `FD1TQHS_TE_CP_SETUP_negedge_posedge, `FD1TQHS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FD1TQHS_TI_CP_SETUP_posedge_posedge, `FD1TQHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FD1TQHS_TI_CP_SETUP_negedge_posedge, `FD1TQHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TEX, posedge D, `FD1TQHS_D_CP_SETUP_posedge_posedge, `FD1TQHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TEX, negedge D, `FD1TQHS_D_CP_SETUP_negedge_posedge, `FD1TQHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD1TQHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1TQHS_CP_PWH, 0, Notifier);
`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FD1TQHS_CP_R_Q_R, `FD1TQHS_CP_R_Q_F);
      (posedge CP => (SO +: Mux21DTITE_)) = (`FD1TQHS_CP_R_SO_R, `FD1TQHS_CP_R_SO_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `FD1TQHS_TE_CP_SETUP_posedge_posedge,`FD1TQHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `FD1TQHS_TE_CP_SETUP_negedge_posedge,`FD1TQHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD1TQHS_TI_CP_SETUP_posedge_posedge, `FD1TQHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD1TQHS_TI_CP_SETUP_negedge_posedge, `FD1TQHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `FD1TQHS_D_CP_SETUP_posedge_posedge, `FD1TQHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `FD1TQHS_D_CP_SETUP_negedge_posedge, `FD1TQHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD1TQHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1TQHS_CP_PWH, 0, Notifier);
 
`endif
   endspecify
`endif


endmodule // FD1TQHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:16 and Version :1.1 //
 
//  START 
// CELL FD1TQHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD1TQHSP_CP_R_SO_R 0.1
`define FD1TQHSP_CP_R_SO_F 0.1
`define FD1TQHSP_CP_R_Q_R 0.1
`define FD1TQHSP_CP_R_Q_F 0.1
`define FD1TQHSP_CP_PWH 0.1
`define FD1TQHSP_CP_PWL 0.1
`define FD1TQHSP_D_CP_SETUP_posedge_posedge 0.1
`define FD1TQHSP_D_CP_SETUP_negedge_posedge 0.1
`define FD1TQHSP_D_CP_HOLD_posedge_posedge 0.1
`define FD1TQHSP_D_CP_HOLD_negedge_posedge 0.1
`define FD1TQHSP_TI_CP_SETUP_posedge_posedge 0.1
`define FD1TQHSP_TI_CP_SETUP_negedge_posedge 0.1
`define FD1TQHSP_TI_CP_HOLD_posedge_posedge 0.1
`define FD1TQHSP_TI_CP_HOLD_negedge_posedge 0.1
`define FD1TQHSP_TE_CP_SETUP_posedge_posedge 0.1
`define FD1TQHSP_TE_CP_SETUP_negedge_posedge 0.1
`define FD1TQHSP_TE_CP_HOLD_posedge_posedge 0.1
`define FD1TQHSP_TE_CP_HOLD_negedge_posedge 0.1

module FD1TQHSP (Q, SO, D, CP, TI, TE);

   output Q;
   output SO;
   input D;
   input CP;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, Notifier);

   buf  u2 (Q, IQ);
buf  u3 (SO, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault

      if(!TE) (posedge CP => (Q +: D)) = (`FD1TQHSP_CP_R_Q_R, `FD1TQHSP_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD1TQHSP_CP_R_Q_R, `FD1TQHSP_CP_R_Q_F);
      if(!D && TI) (posedge CP => (Q +: TE)) = (`FD1TQHSP_CP_R_Q_R, `FD1TQHSP_CP_R_Q_F);
      if(!TI && D) (posedge CP => (Q -: TE)) = (`FD1TQHSP_CP_R_Q_R, `FD1TQHSP_CP_R_Q_F);
      if(!TE) (posedge CP => (SO +: D)) = (`FD1TQHSP_CP_R_SO_R, `FD1TQHSP_CP_R_SO_F);
      if(TE) (posedge CP => (SO +: TI)) = (`FD1TQHSP_CP_R_SO_R, `FD1TQHSP_CP_R_SO_F);
      if(!D && TI) (posedge CP => (SO +: TE)) = (`FD1TQHSP_CP_R_SO_R, `FD1TQHSP_CP_R_SO_F);
      if(!TI && D) (posedge CP => (SO -: TE)) = (`FD1TQHSP_CP_R_SO_R, `FD1TQHSP_CP_R_SO_F);

	$setuphold(posedge CP &&& XorDTI_, posedge TE, `FD1TQHSP_TE_CP_SETUP_posedge_posedge, `FD1TQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& XorDTI_, negedge TE, `FD1TQHSP_TE_CP_SETUP_negedge_posedge, `FD1TQHSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FD1TQHSP_TI_CP_SETUP_posedge_posedge, `FD1TQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FD1TQHSP_TI_CP_SETUP_negedge_posedge, `FD1TQHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TEX, posedge D, `FD1TQHSP_D_CP_SETUP_posedge_posedge, `FD1TQHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TEX, negedge D, `FD1TQHSP_D_CP_SETUP_negedge_posedge, `FD1TQHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD1TQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1TQHSP_CP_PWH, 0, Notifier);
`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FD1TQHSP_CP_R_Q_R, `FD1TQHSP_CP_R_Q_F);
      (posedge CP => (SO +: Mux21DTITE_)) = (`FD1TQHSP_CP_R_SO_R, `FD1TQHSP_CP_R_SO_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `FD1TQHSP_TE_CP_SETUP_posedge_posedge,`FD1TQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `FD1TQHSP_TE_CP_SETUP_negedge_posedge,`FD1TQHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD1TQHSP_TI_CP_SETUP_posedge_posedge, `FD1TQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD1TQHSP_TI_CP_SETUP_negedge_posedge, `FD1TQHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `FD1TQHSP_D_CP_SETUP_posedge_posedge, `FD1TQHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `FD1TQHSP_D_CP_SETUP_negedge_posedge, `FD1TQHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD1TQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1TQHSP_CP_PWH, 0, Notifier);
 
`endif
   endspecify
`endif


endmodule // FD1TQHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:16 and Version :1.1 //
 
//  START 
// CELL FD1TQHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD1TQHSX4_CP_R_SO_R 0.1
`define FD1TQHSX4_CP_R_SO_F 0.1
`define FD1TQHSX4_CP_R_Q_R 0.1
`define FD1TQHSX4_CP_R_Q_F 0.1
`define FD1TQHSX4_CP_PWH 0.1
`define FD1TQHSX4_CP_PWL 0.1
`define FD1TQHSX4_D_CP_SETUP_posedge_posedge 0.1
`define FD1TQHSX4_D_CP_SETUP_negedge_posedge 0.1
`define FD1TQHSX4_D_CP_HOLD_posedge_posedge 0.1
`define FD1TQHSX4_D_CP_HOLD_negedge_posedge 0.1
`define FD1TQHSX4_TI_CP_SETUP_posedge_posedge 0.1
`define FD1TQHSX4_TI_CP_SETUP_negedge_posedge 0.1
`define FD1TQHSX4_TI_CP_HOLD_posedge_posedge 0.1
`define FD1TQHSX4_TI_CP_HOLD_negedge_posedge 0.1
`define FD1TQHSX4_TE_CP_SETUP_posedge_posedge 0.1
`define FD1TQHSX4_TE_CP_SETUP_negedge_posedge 0.1
`define FD1TQHSX4_TE_CP_HOLD_posedge_posedge 0.1
`define FD1TQHSX4_TE_CP_HOLD_negedge_posedge 0.1

module FD1TQHSX4 (Q, SO, D, CP, TI, TE);

   output Q;
   output SO;
   input D;
   input CP;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, Notifier);

   buf  u2 (Q, IQ);
buf  u3 (SO, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault

      if(!TE) (posedge CP => (Q +: D)) = (`FD1TQHSX4_CP_R_Q_R, `FD1TQHSX4_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD1TQHSX4_CP_R_Q_R, `FD1TQHSX4_CP_R_Q_F);
      if(!D && TI) (posedge CP => (Q +: TE)) = (`FD1TQHSX4_CP_R_Q_R, `FD1TQHSX4_CP_R_Q_F);
      if(!TI && D) (posedge CP => (Q -: TE)) = (`FD1TQHSX4_CP_R_Q_R, `FD1TQHSX4_CP_R_Q_F);
      if(!TE) (posedge CP => (SO +: D)) = (`FD1TQHSX4_CP_R_SO_R, `FD1TQHSX4_CP_R_SO_F);
      if(TE) (posedge CP => (SO +: TI)) = (`FD1TQHSX4_CP_R_SO_R, `FD1TQHSX4_CP_R_SO_F);
      if(!D && TI) (posedge CP => (SO +: TE)) = (`FD1TQHSX4_CP_R_SO_R, `FD1TQHSX4_CP_R_SO_F);
      if(!TI && D) (posedge CP => (SO -: TE)) = (`FD1TQHSX4_CP_R_SO_R, `FD1TQHSX4_CP_R_SO_F);

	$setuphold(posedge CP &&& XorDTI_, posedge TE, `FD1TQHSX4_TE_CP_SETUP_posedge_posedge, `FD1TQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& XorDTI_, negedge TE, `FD1TQHSX4_TE_CP_SETUP_negedge_posedge, `FD1TQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FD1TQHSX4_TI_CP_SETUP_posedge_posedge, `FD1TQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FD1TQHSX4_TI_CP_SETUP_negedge_posedge, `FD1TQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TEX, posedge D, `FD1TQHSX4_D_CP_SETUP_posedge_posedge, `FD1TQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TEX, negedge D, `FD1TQHSX4_D_CP_SETUP_negedge_posedge, `FD1TQHSX4_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD1TQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1TQHSX4_CP_PWH, 0, Notifier);
`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FD1TQHSX4_CP_R_Q_R, `FD1TQHSX4_CP_R_Q_F);
      (posedge CP => (SO +: Mux21DTITE_)) = (`FD1TQHSX4_CP_R_SO_R, `FD1TQHSX4_CP_R_SO_F);
 
        $setuphold(posedge CP &&& XorDTI_, posedge TE, `FD1TQHSX4_TE_CP_SETUP_posedge_posedge,`FD1TQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& XorDTI_, negedge TE, `FD1TQHSX4_TE_CP_SETUP_negedge_posedge,`FD1TQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD1TQHSX4_TI_CP_SETUP_posedge_posedge, `FD1TQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD1TQHSX4_TI_CP_SETUP_negedge_posedge, `FD1TQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge D, `FD1TQHSX4_D_CP_SETUP_posedge_posedge, `FD1TQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge D, `FD1TQHSX4_D_CP_SETUP_negedge_posedge, `FD1TQHSX4_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD1TQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD1TQHSX4_CP_PWH, 0, Notifier);
 
`endif
   endspecify
`endif


endmodule // FD1TQHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:16 and Version :1.1 //
 
//  START 
// CELL FD2HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD2HS_CD_F_QN_R 0.1
`define FD2HS_CP_R_QN_F 0.1
`define FD2HS_CP_R_QN_R 0.1
`define FD2HS_CD_F_Q_F 0.1
`define FD2HS_CP_R_Q_R 0.1
`define FD2HS_CP_R_Q_F 0.1
`define FD2HS_CD_CP_REM_posedge_posedge 0.1
`define FD2HS_CD_CP_REC_posedge_posedge 0.1
`define FD2HS_CD_PWL 0.1
`define FD2HS_CP_PWH 0.1
`define FD2HS_CP_PWL 0.1
`define FD2HS_D_CP_SETUP_posedge_posedge 0.1
`define FD2HS_D_CP_SETUP_negedge_posedge 0.1
`define FD2HS_D_CP_HOLD_posedge_posedge 0.1
`define FD2HS_D_CP_HOLD_negedge_posedge 0.1

module FD2HS (Q, QN, D, CP, CD);

   output Q;
   output QN;
   input D;
   input CP;
   input CD;


   reg Notifier;


   U_FD_P_RN_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, CD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(CD) (posedge CP => (Q +: D)) = (`FD2HS_CP_R_Q_R, `FD2HS_CP_R_Q_F);
      if(CD) (posedge CP => (QN -: D)) = (`FD2HS_CP_R_QN_R, `FD2HS_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2HS_CD_F_Q_F,`FD2HS_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FD2HS_CD_F_QN_R,`FD2HS_CD_F_QN_R);

	$setuphold(posedge CP &&& CD, posedge D, `FD2HS_D_CP_SETUP_posedge_posedge, `FD2HS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge D, `FD2HS_D_CP_SETUP_negedge_posedge, `FD2HS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD2HS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2HS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2HS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& D, `FD2HS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D, posedge CD, `FD2HS_CD_CP_REM_posedge_posedge, Notifier);
`else

      (posedge CP => (Q +: D)) = (`FD2HS_CP_R_Q_R, `FD2HS_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`FD2HS_CP_R_QN_R, `FD2HS_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2HS_CD_F_Q_F,`FD2HS_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FD2HS_CD_F_QN_R,`FD2HS_CD_F_QN_R);
 
        $setuphold(posedge CP &&& CD, posedge D, `FD2HS_D_CP_SETUP_posedge_posedge, `FD2HS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge D, `FD2HS_D_CP_SETUP_negedge_posedge, `FD2HS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD2HS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2HS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2HS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& D, `FD2HS_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D, posedge CD, `FD2HS_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FD2HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:20 and Version :1.1 //
 
//  START 
// CELL FD2HSP

`celldefine
// `define functional //off sdf
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD2HSP_CD_F_QN_R 0.1
`define FD2HSP_CP_R_QN_F 0.1
`define FD2HSP_CP_R_QN_R 0.1
`define FD2HSP_CD_F_Q_F 0.1
`define FD2HSP_CP_R_Q_R 0.1
`define FD2HSP_CP_R_Q_F 0.1
`define FD2HSP_CD_CP_REM_posedge_posedge 0.1
`define FD2HSP_CD_CP_REC_posedge_posedge 0.1
`define FD2HSP_CD_PWL 0.1
`define FD2HSP_CP_PWH 0.1
`define FD2HSP_CP_PWL 0.1
`define FD2HSP_D_CP_SETUP_posedge_posedge 0.1
`define FD2HSP_D_CP_SETUP_negedge_posedge 0.1
`define FD2HSP_D_CP_HOLD_posedge_posedge 0.1
`define FD2HSP_D_CP_HOLD_negedge_posedge 0.1

module FD2HSP (Q, QN, D, CP, CD);

   output Q;
   output QN;
   input D;
   input CP;
   input CD;


   reg Notifier;


   U_FD_P_RN_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, CD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(CD) (posedge CP => (Q +: D)) = (`FD2HSP_CP_R_Q_R, `FD2HSP_CP_R_Q_F);
      if(CD) (posedge CP => (QN -: D)) = (`FD2HSP_CP_R_QN_R, `FD2HSP_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2HSP_CD_F_Q_F,`FD2HSP_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FD2HSP_CD_F_QN_R,`FD2HSP_CD_F_QN_R);

	// $setuphold(posedge CP &&& CD, posedge D, `FD2HSP_D_CP_SETUP_posedge_posedge, `FD2HSP_D_CP_HOLD_posedge_posedge, Notifier);
	// $setuphold(posedge CP &&& CD, negedge D, `FD2HSP_D_CP_SETUP_negedge_posedge, `FD2HSP_D_CP_HOLD_negedge_posedge, Notifier);

   //    $width(negedge CP, `FD2HSP_CP_PWL, 0, Notifier);
   //    $width(posedge CP &&& CD, `FD2HSP_CP_PWH, 0, Notifier);
   //    $width(negedge CD, `FD2HSP_CD_PWL, 0, Notifier);
	// $recovery(posedge CD, posedge CP &&& D, `FD2HSP_CD_CP_REC_posedge_posedge, Notifier);

	// $hold(posedge CP &&& D, posedge CD, `FD2HSP_CD_CP_REM_posedge_posedge, Notifier);
`else

      (posedge CP => (Q +: D)) = (`FD2HSP_CP_R_Q_R, `FD2HSP_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`FD2HSP_CP_R_QN_R, `FD2HSP_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2HSP_CD_F_Q_F,`FD2HSP_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FD2HSP_CD_F_QN_R,`FD2HSP_CD_F_QN_R);
 
      //   $setuphold(posedge CP &&& CD, posedge D, `FD2HSP_D_CP_SETUP_posedge_posedge, `FD2HSP_D_CP_HOLD_posedge_posedge, Notifier);
      //   $setuphold(posedge CP &&& CD, negedge D, `FD2HSP_D_CP_SETUP_negedge_posedge, `FD2HSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      // $width(negedge CP, `FD2HSP_CP_PWL, 0, Notifier);
      // $width(posedge CP &&& CD, `FD2HSP_CP_PWH, 0, Notifier);
      // $width(negedge CD, `FD2HSP_CD_PWL, 0, Notifier);
      //   $recovery(posedge CD, posedge CP &&& D, `FD2HSP_CD_CP_REC_posedge_posedge, Notifier);
 
      //   $hold(posedge CP &&& D, posedge CD, `FD2HSP_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FD2HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:20 and Version :1.1 //
 
//  START 
// CELL FDM2HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDM2HS_CD_F_QN_R 0.1
`define FDM2HS_CP_R_QN_F 0.1
`define FDM2HS_CP_R_QN_R 0.1
`define FDM2HS_CD_F_Q_F 0.1
`define FDM2HS_CP_R_Q_R 0.1
`define FDM2HS_CP_R_Q_F 0.1
`define FDM2HS_CD_CP_REM_posedge_posedge 0.1
`define FDM2HS_CD_CP_REC_posedge_posedge 0.1
`define FDM2HS_CD_PWL 0.1
`define FDM2HS_CP_PWH 0.1
`define FDM2HS_CP_PWL 0.1
`define FDM2HS_D_CP_SETUP_posedge_posedge 0.1
`define FDM2HS_D_CP_SETUP_negedge_posedge 0.1
`define FDM2HS_D_CP_HOLD_posedge_posedge 0.1
`define FDM2HS_D_CP_HOLD_negedge_posedge 0.1

module FDM2HS (Q, QN, D, CP, CD);

   output Q;
   output QN;
   input D;
   input CP;
   input CD;


   reg Notifier;


   U_FD_P_RN_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, CD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(CD) (posedge CP => (Q +: D)) = (`FDM2HS_CP_R_Q_R, `FDM2HS_CP_R_Q_F);
      if(CD) (posedge CP => (QN -: D)) = (`FDM2HS_CP_R_QN_R, `FDM2HS_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FDM2HS_CD_F_Q_F,`FDM2HS_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FDM2HS_CD_F_QN_R,`FDM2HS_CD_F_QN_R);

	$setuphold(posedge CP &&& CD, posedge D, `FDM2HS_D_CP_SETUP_posedge_posedge, `FDM2HS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge D, `FDM2HS_D_CP_SETUP_negedge_posedge, `FDM2HS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDM2HS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDM2HS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDM2HS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& D, `FDM2HS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D, posedge CD, `FDM2HS_CD_CP_REM_posedge_posedge, Notifier);
`else

      (posedge CP => (Q +: D)) = (`FDM2HS_CP_R_Q_R, `FDM2HS_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`FDM2HS_CP_R_QN_R, `FDM2HS_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FDM2HS_CD_F_Q_F,`FDM2HS_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FDM2HS_CD_F_QN_R,`FDM2HS_CD_F_QN_R);
 
        $setuphold(posedge CP &&& CD, posedge D, `FDM2HS_D_CP_SETUP_posedge_posedge, `FDM2HS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge D, `FDM2HS_D_CP_SETUP_negedge_posedge, `FDM2HS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDM2HS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDM2HS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDM2HS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& D, `FDM2HS_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D, posedge CD, `FDM2HS_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FDM2HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:20 and Version :1.1 //
 
//  START 
// CELL FDM2HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDM2HSP_CD_F_QN_R 0.1
`define FDM2HSP_CP_R_QN_F 0.1
`define FDM2HSP_CP_R_QN_R 0.1
`define FDM2HSP_CD_F_Q_F 0.1
`define FDM2HSP_CP_R_Q_R 0.1
`define FDM2HSP_CP_R_Q_F 0.1
`define FDM2HSP_CD_CP_REM_posedge_posedge 0.1
`define FDM2HSP_CD_CP_REC_posedge_posedge 0.1
`define FDM2HSP_CD_PWL 0.1
`define FDM2HSP_CP_PWH 0.1
`define FDM2HSP_CP_PWL 0.1
`define FDM2HSP_D_CP_SETUP_posedge_posedge 0.1
`define FDM2HSP_D_CP_SETUP_negedge_posedge 0.1
`define FDM2HSP_D_CP_HOLD_posedge_posedge 0.1
`define FDM2HSP_D_CP_HOLD_negedge_posedge 0.1

module FDM2HSP (Q, QN, D, CP, CD);

   output Q;
   output QN;
   input D;
   input CP;
   input CD;


   reg Notifier;


   U_FD_P_RN_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, CD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(CD) (posedge CP => (Q +: D)) = (`FDM2HSP_CP_R_Q_R, `FDM2HSP_CP_R_Q_F);
      if(CD) (posedge CP => (QN -: D)) = (`FDM2HSP_CP_R_QN_R, `FDM2HSP_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FDM2HSP_CD_F_Q_F,`FDM2HSP_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FDM2HSP_CD_F_QN_R,`FDM2HSP_CD_F_QN_R);

	$setuphold(posedge CP &&& CD, posedge D, `FDM2HSP_D_CP_SETUP_posedge_posedge, `FDM2HSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge D, `FDM2HSP_D_CP_SETUP_negedge_posedge, `FDM2HSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDM2HSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDM2HSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDM2HSP_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& D, `FDM2HSP_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D, posedge CD, `FDM2HSP_CD_CP_REM_posedge_posedge, Notifier);
`else

      (posedge CP => (Q +: D)) = (`FDM2HSP_CP_R_Q_R, `FDM2HSP_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`FDM2HSP_CP_R_QN_R, `FDM2HSP_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FDM2HSP_CD_F_Q_F,`FDM2HSP_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FDM2HSP_CD_F_QN_R,`FDM2HSP_CD_F_QN_R);
 
        $setuphold(posedge CP &&& CD, posedge D, `FDM2HSP_D_CP_SETUP_posedge_posedge, `FDM2HSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge D, `FDM2HSP_D_CP_SETUP_negedge_posedge, `FDM2HSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDM2HSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDM2HSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDM2HSP_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& D, `FDM2HSP_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D, posedge CD, `FDM2HSP_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FDM2HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:20 and Version :1.1 //
 
//  START 
// CELL FDH2HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDH2HSX4_CD_F_QN_R 0.1
`define FDH2HSX4_CP_R_QN_F 0.1
`define FDH2HSX4_CP_R_QN_R 0.1
`define FDH2HSX4_CD_F_Q_F 0.1
`define FDH2HSX4_CP_R_Q_R 0.1
`define FDH2HSX4_CP_R_Q_F 0.1
`define FDH2HSX4_CD_CP_REM_posedge_posedge 0.1
`define FDH2HSX4_CD_CP_REC_posedge_posedge 0.1
`define FDH2HSX4_CD_PWL 0.1
`define FDH2HSX4_CP_PWH 0.1
`define FDH2HSX4_CP_PWL 0.1
`define FDH2HSX4_D_CP_SETUP_posedge_posedge 0.1
`define FDH2HSX4_D_CP_SETUP_negedge_posedge 0.1
`define FDH2HSX4_D_CP_HOLD_posedge_posedge 0.1
`define FDH2HSX4_D_CP_HOLD_negedge_posedge 0.1

module FDH2HSX4 (Q, QN, D, CP, CD);

   output Q;
   output QN;
   input D;
   input CP;
   input CD;


   reg Notifier;


   U_FD_P_RN_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, CD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(CD) (posedge CP => (Q +: D)) = (`FDH2HSX4_CP_R_Q_R, `FDH2HSX4_CP_R_Q_F);
      if(CD) (posedge CP => (QN -: D)) = (`FDH2HSX4_CP_R_QN_R, `FDH2HSX4_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FDH2HSX4_CD_F_Q_F,`FDH2HSX4_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FDH2HSX4_CD_F_QN_R,`FDH2HSX4_CD_F_QN_R);

	$setuphold(posedge CP &&& CD, posedge D, `FDH2HSX4_D_CP_SETUP_posedge_posedge, `FDH2HSX4_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge D, `FDH2HSX4_D_CP_SETUP_negedge_posedge, `FDH2HSX4_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDH2HSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDH2HSX4_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDH2HSX4_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& D, `FDH2HSX4_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D, posedge CD, `FDH2HSX4_CD_CP_REM_posedge_posedge, Notifier);
`else

      (posedge CP => (Q +: D)) = (`FDH2HSX4_CP_R_Q_R, `FDH2HSX4_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`FDH2HSX4_CP_R_QN_R, `FDH2HSX4_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FDH2HSX4_CD_F_Q_F,`FDH2HSX4_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FDH2HSX4_CD_F_QN_R,`FDH2HSX4_CD_F_QN_R);
 
        $setuphold(posedge CP &&& CD, posedge D, `FDH2HSX4_D_CP_SETUP_posedge_posedge, `FDH2HSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge D, `FDH2HSX4_D_CP_SETUP_negedge_posedge, `FDH2HSX4_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDH2HSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDH2HSX4_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDH2HSX4_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& D, `FDH2HSX4_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D, posedge CD, `FDH2HSX4_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FDH2HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:20 and Version :1.1 //
 
//  START 
// CELL FDH2HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDH2HSX8_CD_F_QN_R 0.1
`define FDH2HSX8_CP_R_QN_F 0.1
`define FDH2HSX8_CP_R_QN_R 0.1
`define FDH2HSX8_CD_F_Q_F 0.1
`define FDH2HSX8_CP_R_Q_R 0.1
`define FDH2HSX8_CP_R_Q_F 0.1
`define FDH2HSX8_CD_CP_REM_posedge_posedge 0.1
`define FDH2HSX8_CD_CP_REC_posedge_posedge 0.1
`define FDH2HSX8_CD_PWL 0.1
`define FDH2HSX8_CP_PWH 0.1
`define FDH2HSX8_CP_PWL 0.1
`define FDH2HSX8_D_CP_SETUP_posedge_posedge 0.1
`define FDH2HSX8_D_CP_SETUP_negedge_posedge 0.1
`define FDH2HSX8_D_CP_HOLD_posedge_posedge 0.1
`define FDH2HSX8_D_CP_HOLD_negedge_posedge 0.1

module FDH2HSX8 (Q, QN, D, CP, CD);

   output Q;
   output QN;
   input D;
   input CP;
   input CD;


   reg Notifier;


   U_FD_P_RN_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, CD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(CD) (posedge CP => (Q +: D)) = (`FDH2HSX8_CP_R_Q_R, `FDH2HSX8_CP_R_Q_F);
      if(CD) (posedge CP => (QN -: D)) = (`FDH2HSX8_CP_R_QN_R, `FDH2HSX8_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FDH2HSX8_CD_F_Q_F,`FDH2HSX8_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FDH2HSX8_CD_F_QN_R,`FDH2HSX8_CD_F_QN_R);

	$setuphold(posedge CP &&& CD, posedge D, `FDH2HSX8_D_CP_SETUP_posedge_posedge, `FDH2HSX8_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge D, `FDH2HSX8_D_CP_SETUP_negedge_posedge, `FDH2HSX8_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDH2HSX8_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDH2HSX8_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDH2HSX8_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& D, `FDH2HSX8_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D, posedge CD, `FDH2HSX8_CD_CP_REM_posedge_posedge, Notifier);
`else

      (posedge CP => (Q +: D)) = (`FDH2HSX8_CP_R_Q_R, `FDH2HSX8_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`FDH2HSX8_CP_R_QN_R, `FDH2HSX8_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FDH2HSX8_CD_F_Q_F,`FDH2HSX8_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FDH2HSX8_CD_F_QN_R,`FDH2HSX8_CD_F_QN_R);
 
        $setuphold(posedge CP &&& CD, posedge D, `FDH2HSX8_D_CP_SETUP_posedge_posedge, `FDH2HSX8_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge D, `FDH2HSX8_D_CP_SETUP_negedge_posedge, `FDH2HSX8_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDH2HSX8_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDH2HSX8_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDH2HSX8_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& D, `FDH2HSX8_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D, posedge CD, `FDH2HSX8_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FDH2HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:20 and Version :1.1 //
 
//  START 
// CELL F_FD2HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_FD2HS_CD_F_QN_R 0.1
`define F_FD2HS_CP_R_QN_F 0.1
`define F_FD2HS_CP_R_QN_R 0.1
`define F_FD2HS_CD_F_Q_F 0.1
`define F_FD2HS_CP_R_Q_R 0.1
`define F_FD2HS_CP_R_Q_F 0.1
`define F_FD2HS_CD_CP_REM_posedge_posedge 0.1
`define F_FD2HS_CD_CP_REC_posedge_posedge 0.1
`define F_FD2HS_CD_PWL 0.1
`define F_FD2HS_CP_PWH 0.1
`define F_FD2HS_CP_PWL 0.1
`define F_FD2HS_D_CP_SETUP_posedge_posedge 0.1
`define F_FD2HS_D_CP_SETUP_negedge_posedge 0.1
`define F_FD2HS_D_CP_HOLD_posedge_posedge 0.1
`define F_FD2HS_D_CP_HOLD_negedge_posedge 0.1

module F_FD2HS (Q, QN, D, CP, CD);

   output Q;
   output QN;
   input D;
   input CP;
   input CD;


   reg Notifier;


   U_FD_P_RN_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, CD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(CD) (posedge CP => (Q +: D)) = (`F_FD2HS_CP_R_Q_R, `F_FD2HS_CP_R_Q_F);
      if(CD) (posedge CP => (QN -: D)) = (`F_FD2HS_CP_R_QN_R, `F_FD2HS_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`F_FD2HS_CD_F_Q_F,`F_FD2HS_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`F_FD2HS_CD_F_QN_R,`F_FD2HS_CD_F_QN_R);

	$setuphold(posedge CP &&& CD, posedge D, `F_FD2HS_D_CP_SETUP_posedge_posedge, `F_FD2HS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge D, `F_FD2HS_D_CP_SETUP_negedge_posedge, `F_FD2HS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `F_FD2HS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `F_FD2HS_CP_PWH, 0, Notifier);
      $width(negedge CD, `F_FD2HS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& D, `F_FD2HS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D, posedge CD, `F_FD2HS_CD_CP_REM_posedge_posedge, Notifier);
`else

      (posedge CP => (Q +: D)) = (`F_FD2HS_CP_R_Q_R, `F_FD2HS_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`F_FD2HS_CP_R_QN_R, `F_FD2HS_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`F_FD2HS_CD_F_Q_F,`F_FD2HS_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`F_FD2HS_CD_F_QN_R,`F_FD2HS_CD_F_QN_R);
 
        $setuphold(posedge CP &&& CD, posedge D, `F_FD2HS_D_CP_SETUP_posedge_posedge, `F_FD2HS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge D, `F_FD2HS_D_CP_SETUP_negedge_posedge, `F_FD2HS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `F_FD2HS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `F_FD2HS_CP_PWH, 0, Notifier);
      $width(negedge CD, `F_FD2HS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& D, `F_FD2HS_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D, posedge CD, `F_FD2HS_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // F_FD2HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:20 and Version :1.1 //
 
//  START 
// CELL F_FD2HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_FD2HSP_CD_F_QN_R 0.1
`define F_FD2HSP_CP_R_QN_F 0.1
`define F_FD2HSP_CP_R_QN_R 0.1
`define F_FD2HSP_CD_F_Q_F 0.1
`define F_FD2HSP_CP_R_Q_R 0.1
`define F_FD2HSP_CP_R_Q_F 0.1
`define F_FD2HSP_CD_CP_REM_posedge_posedge 0.1
`define F_FD2HSP_CD_CP_REC_posedge_posedge 0.1
`define F_FD2HSP_CD_PWL 0.1
`define F_FD2HSP_CP_PWH 0.1
`define F_FD2HSP_CP_PWL 0.1
`define F_FD2HSP_D_CP_SETUP_posedge_posedge 0.1
`define F_FD2HSP_D_CP_SETUP_negedge_posedge 0.1
`define F_FD2HSP_D_CP_HOLD_posedge_posedge 0.1
`define F_FD2HSP_D_CP_HOLD_negedge_posedge 0.1

module F_FD2HSP (Q, QN, D, CP, CD);

   output Q;
   output QN;
   input D;
   input CP;
   input CD;


   reg Notifier;


   U_FD_P_RN_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, CD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(CD) (posedge CP => (Q +: D)) = (`F_FD2HSP_CP_R_Q_R, `F_FD2HSP_CP_R_Q_F);
      if(CD) (posedge CP => (QN -: D)) = (`F_FD2HSP_CP_R_QN_R, `F_FD2HSP_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`F_FD2HSP_CD_F_Q_F,`F_FD2HSP_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`F_FD2HSP_CD_F_QN_R,`F_FD2HSP_CD_F_QN_R);

	$setuphold(posedge CP &&& CD, posedge D, `F_FD2HSP_D_CP_SETUP_posedge_posedge, `F_FD2HSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge D, `F_FD2HSP_D_CP_SETUP_negedge_posedge, `F_FD2HSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `F_FD2HSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `F_FD2HSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `F_FD2HSP_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& D, `F_FD2HSP_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D, posedge CD, `F_FD2HSP_CD_CP_REM_posedge_posedge, Notifier);
`else

      (posedge CP => (Q +: D)) = (`F_FD2HSP_CP_R_Q_R, `F_FD2HSP_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`F_FD2HSP_CP_R_QN_R, `F_FD2HSP_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`F_FD2HSP_CD_F_Q_F,`F_FD2HSP_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`F_FD2HSP_CD_F_QN_R,`F_FD2HSP_CD_F_QN_R);
 
        $setuphold(posedge CP &&& CD, posedge D, `F_FD2HSP_D_CP_SETUP_posedge_posedge, `F_FD2HSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge D, `F_FD2HSP_D_CP_SETUP_negedge_posedge, `F_FD2HSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `F_FD2HSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `F_FD2HSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `F_FD2HSP_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& D, `F_FD2HSP_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D, posedge CD, `F_FD2HSP_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // F_FD2HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:20 and Version :1.1 //
 
//  START 
// CELL FD2QHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD2QHS_CD_F_Q_F 0.1
`define FD2QHS_CP_R_Q_R 0.1
`define FD2QHS_CP_R_Q_F 0.1
`define FD2QHS_D_CP_HOLD_posedge_posedge 0.1
`define FD2QHS_D_CP_HOLD_negedge_posedge 0.1
`define FD2QHS_D_CP_SETUP_posedge_posedge 0.1
`define FD2QHS_D_CP_SETUP_negedge_posedge 0.1
`define FD2QHS_CP_PWL 0.1
`define FD2QHS_CP_PWH 0.1
`define FD2QHS_CD_PWL 0.1
`define FD2QHS_CD_CP_REC_posedge_posedge 0.1
`define FD2QHS_CD_CP_REM_posedge_posedge 0.1

module FD2QHS (Q, D, CP, CD);

   output Q;
   input D;
   input CP;
   input CD;


   reg Notifier;


   U_FD_P_RN_NOTI u0 (IQ, D, CP, CD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(CD) (posedge CP => (Q +: D)) = (`FD2QHS_CP_R_Q_R, `FD2QHS_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2QHS_CD_F_Q_F,`FD2QHS_CD_F_Q_F);

	$setuphold(posedge CP &&& CD, posedge D, `FD2QHS_D_CP_SETUP_posedge_posedge, `FD2QHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge D, `FD2QHS_D_CP_SETUP_negedge_posedge, `FD2QHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD2QHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2QHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2QHS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& D, `FD2QHS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D, posedge CD, `FD2QHS_CD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: D)) = (`FD2QHS_CP_R_Q_R, `FD2QHS_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2QHS_CD_F_Q_F,`FD2QHS_CD_F_Q_F);
 
        $setuphold(posedge CP &&& CD, posedge D, `FD2QHS_D_CP_SETUP_posedge_posedge, `FD2QHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge D, `FD2QHS_D_CP_SETUP_negedge_posedge, `FD2QHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD2QHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2QHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2QHS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& D, `FD2QHS_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D, posedge CD, `FD2QHS_CD_CP_REM_posedge_posedge, Notifier);
 
`endif
   endspecify
`endif


endmodule // FD2QHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:27 and Version :1.1 //
 
//  START 
// CELL FD2QHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD2QHSP_CD_F_Q_F 0.1
`define FD2QHSP_CP_R_Q_R 0.1
`define FD2QHSP_CP_R_Q_F 0.1
`define FD2QHSP_D_CP_HOLD_posedge_posedge 0.1
`define FD2QHSP_D_CP_HOLD_negedge_posedge 0.1
`define FD2QHSP_D_CP_SETUP_posedge_posedge 0.1
`define FD2QHSP_D_CP_SETUP_negedge_posedge 0.1
`define FD2QHSP_CP_PWL 0.1
`define FD2QHSP_CP_PWH 0.1
`define FD2QHSP_CD_PWL 0.1
`define FD2QHSP_CD_CP_REC_posedge_posedge 0.1
`define FD2QHSP_CD_CP_REM_posedge_posedge 0.1

module FD2QHSP (Q, D, CP, CD);

   output Q;
   input D;
   input CP;
   input CD;


   reg Notifier;


   U_FD_P_RN_NOTI u0 (IQ, D, CP, CD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(CD) (posedge CP => (Q +: D)) = (`FD2QHSP_CP_R_Q_R, `FD2QHSP_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2QHSP_CD_F_Q_F,`FD2QHSP_CD_F_Q_F);

	$setuphold(posedge CP &&& CD, posedge D, `FD2QHSP_D_CP_SETUP_posedge_posedge, `FD2QHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge D, `FD2QHSP_D_CP_SETUP_negedge_posedge, `FD2QHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD2QHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2QHSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2QHSP_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& D, `FD2QHSP_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D, posedge CD, `FD2QHSP_CD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: D)) = (`FD2QHSP_CP_R_Q_R, `FD2QHSP_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2QHSP_CD_F_Q_F,`FD2QHSP_CD_F_Q_F);
 
        $setuphold(posedge CP &&& CD, posedge D, `FD2QHSP_D_CP_SETUP_posedge_posedge, `FD2QHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge D, `FD2QHSP_D_CP_SETUP_negedge_posedge, `FD2QHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD2QHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2QHSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2QHSP_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& D, `FD2QHSP_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D, posedge CD, `FD2QHSP_CD_CP_REM_posedge_posedge, Notifier);
 
`endif
   endspecify
`endif


endmodule // FD2QHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:27 and Version :1.1 //
 
//  START 
// CELL FD2QHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD2QHSX4_CD_F_Q_F 0.1
`define FD2QHSX4_CP_R_Q_R 0.1
`define FD2QHSX4_CP_R_Q_F 0.1
`define FD2QHSX4_D_CP_HOLD_posedge_posedge 0.1
`define FD2QHSX4_D_CP_HOLD_negedge_posedge 0.1
`define FD2QHSX4_D_CP_SETUP_posedge_posedge 0.1
`define FD2QHSX4_D_CP_SETUP_negedge_posedge 0.1
`define FD2QHSX4_CP_PWL 0.1
`define FD2QHSX4_CP_PWH 0.1
`define FD2QHSX4_CD_PWL 0.1
`define FD2QHSX4_CD_CP_REC_posedge_posedge 0.1
`define FD2QHSX4_CD_CP_REM_posedge_posedge 0.1

module FD2QHSX4 (Q, D, CP, CD);

   output Q;
   input D;
   input CP;
   input CD;


   reg Notifier;


   U_FD_P_RN_NOTI u0 (IQ, D, CP, CD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(CD) (posedge CP => (Q +: D)) = (`FD2QHSX4_CP_R_Q_R, `FD2QHSX4_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2QHSX4_CD_F_Q_F,`FD2QHSX4_CD_F_Q_F);

	$setuphold(posedge CP &&& CD, posedge D, `FD2QHSX4_D_CP_SETUP_posedge_posedge, `FD2QHSX4_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge D, `FD2QHSX4_D_CP_SETUP_negedge_posedge, `FD2QHSX4_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD2QHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2QHSX4_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2QHSX4_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& D, `FD2QHSX4_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D, posedge CD, `FD2QHSX4_CD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: D)) = (`FD2QHSX4_CP_R_Q_R, `FD2QHSX4_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2QHSX4_CD_F_Q_F,`FD2QHSX4_CD_F_Q_F);
 
        $setuphold(posedge CP &&& CD, posedge D, `FD2QHSX4_D_CP_SETUP_posedge_posedge, `FD2QHSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge D, `FD2QHSX4_D_CP_SETUP_negedge_posedge, `FD2QHSX4_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD2QHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2QHSX4_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2QHSX4_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& D, `FD2QHSX4_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D, posedge CD, `FD2QHSX4_CD_CP_REM_posedge_posedge, Notifier);
 
`endif
   endspecify
`endif


endmodule // FD2QHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:27 and Version :1.1 //
 
//  START 
// CELL FDM2QHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDM2QHS_CD_F_Q_F 0.1
`define FDM2QHS_CP_R_Q_R 0.1
`define FDM2QHS_CP_R_Q_F 0.1
`define FDM2QHS_D_CP_HOLD_posedge_posedge 0.1
`define FDM2QHS_D_CP_HOLD_negedge_posedge 0.1
`define FDM2QHS_D_CP_SETUP_posedge_posedge 0.1
`define FDM2QHS_D_CP_SETUP_negedge_posedge 0.1
`define FDM2QHS_CP_PWL 0.1
`define FDM2QHS_CP_PWH 0.1
`define FDM2QHS_CD_PWL 0.1
`define FDM2QHS_CD_CP_REC_posedge_posedge 0.1
`define FDM2QHS_CD_CP_REM_posedge_posedge 0.1

module FDM2QHS (Q, D, CP, CD);

   output Q;
   input D;
   input CP;
   input CD;


   reg Notifier;


   U_FD_P_RN_NOTI u0 (IQ, D, CP, CD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(CD) (posedge CP => (Q +: D)) = (`FDM2QHS_CP_R_Q_R, `FDM2QHS_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FDM2QHS_CD_F_Q_F,`FDM2QHS_CD_F_Q_F);

	$setuphold(posedge CP &&& CD, posedge D, `FDM2QHS_D_CP_SETUP_posedge_posedge, `FDM2QHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge D, `FDM2QHS_D_CP_SETUP_negedge_posedge, `FDM2QHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDM2QHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDM2QHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDM2QHS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& D, `FDM2QHS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D, posedge CD, `FDM2QHS_CD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: D)) = (`FDM2QHS_CP_R_Q_R, `FDM2QHS_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FDM2QHS_CD_F_Q_F,`FDM2QHS_CD_F_Q_F);
 
        $setuphold(posedge CP &&& CD, posedge D, `FDM2QHS_D_CP_SETUP_posedge_posedge, `FDM2QHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge D, `FDM2QHS_D_CP_SETUP_negedge_posedge, `FDM2QHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDM2QHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDM2QHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDM2QHS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& D, `FDM2QHS_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D, posedge CD, `FDM2QHS_CD_CP_REM_posedge_posedge, Notifier);
 
`endif
   endspecify
`endif


endmodule // FDM2QHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:27 and Version :1.1 //
 
//  START 
// CELL FDM2QHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDM2QHSP_CD_F_Q_F 0.1
`define FDM2QHSP_CP_R_Q_R 0.1
`define FDM2QHSP_CP_R_Q_F 0.1
`define FDM2QHSP_D_CP_HOLD_posedge_posedge 0.1
`define FDM2QHSP_D_CP_HOLD_negedge_posedge 0.1
`define FDM2QHSP_D_CP_SETUP_posedge_posedge 0.1
`define FDM2QHSP_D_CP_SETUP_negedge_posedge 0.1
`define FDM2QHSP_CP_PWL 0.1
`define FDM2QHSP_CP_PWH 0.1
`define FDM2QHSP_CD_PWL 0.1
`define FDM2QHSP_CD_CP_REC_posedge_posedge 0.1
`define FDM2QHSP_CD_CP_REM_posedge_posedge 0.1

module FDM2QHSP (Q, D, CP, CD);

   output Q;
   input D;
   input CP;
   input CD;


   reg Notifier;


   U_FD_P_RN_NOTI u0 (IQ, D, CP, CD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(CD) (posedge CP => (Q +: D)) = (`FDM2QHSP_CP_R_Q_R, `FDM2QHSP_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FDM2QHSP_CD_F_Q_F,`FDM2QHSP_CD_F_Q_F);

	$setuphold(posedge CP &&& CD, posedge D, `FDM2QHSP_D_CP_SETUP_posedge_posedge, `FDM2QHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge D, `FDM2QHSP_D_CP_SETUP_negedge_posedge, `FDM2QHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDM2QHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDM2QHSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDM2QHSP_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& D, `FDM2QHSP_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D, posedge CD, `FDM2QHSP_CD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: D)) = (`FDM2QHSP_CP_R_Q_R, `FDM2QHSP_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FDM2QHSP_CD_F_Q_F,`FDM2QHSP_CD_F_Q_F);
 
        $setuphold(posedge CP &&& CD, posedge D, `FDM2QHSP_D_CP_SETUP_posedge_posedge, `FDM2QHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge D, `FDM2QHSP_D_CP_SETUP_negedge_posedge, `FDM2QHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDM2QHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDM2QHSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDM2QHSP_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& D, `FDM2QHSP_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D, posedge CD, `FDM2QHSP_CD_CP_REM_posedge_posedge, Notifier);
 
`endif
   endspecify
`endif


endmodule // FDM2QHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:27 and Version :1.1 //
 
//  START 
// CELL FDH2QHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDH2QHSX4_CD_F_Q_F 0.1
`define FDH2QHSX4_CP_R_Q_R 0.1
`define FDH2QHSX4_CP_R_Q_F 0.1
`define FDH2QHSX4_D_CP_HOLD_posedge_posedge 0.1
`define FDH2QHSX4_D_CP_HOLD_negedge_posedge 0.1
`define FDH2QHSX4_D_CP_SETUP_posedge_posedge 0.1
`define FDH2QHSX4_D_CP_SETUP_negedge_posedge 0.1
`define FDH2QHSX4_CP_PWL 0.1
`define FDH2QHSX4_CP_PWH 0.1
`define FDH2QHSX4_CD_PWL 0.1
`define FDH2QHSX4_CD_CP_REC_posedge_posedge 0.1
`define FDH2QHSX4_CD_CP_REM_posedge_posedge 0.1

module FDH2QHSX4 (Q, D, CP, CD);

   output Q;
   input D;
   input CP;
   input CD;


   reg Notifier;


   U_FD_P_RN_NOTI u0 (IQ, D, CP, CD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(CD) (posedge CP => (Q +: D)) = (`FDH2QHSX4_CP_R_Q_R, `FDH2QHSX4_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FDH2QHSX4_CD_F_Q_F,`FDH2QHSX4_CD_F_Q_F);

	$setuphold(posedge CP &&& CD, posedge D, `FDH2QHSX4_D_CP_SETUP_posedge_posedge, `FDH2QHSX4_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge D, `FDH2QHSX4_D_CP_SETUP_negedge_posedge, `FDH2QHSX4_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDH2QHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDH2QHSX4_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDH2QHSX4_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& D, `FDH2QHSX4_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D, posedge CD, `FDH2QHSX4_CD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: D)) = (`FDH2QHSX4_CP_R_Q_R, `FDH2QHSX4_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FDH2QHSX4_CD_F_Q_F,`FDH2QHSX4_CD_F_Q_F);
 
        $setuphold(posedge CP &&& CD, posedge D, `FDH2QHSX4_D_CP_SETUP_posedge_posedge, `FDH2QHSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge D, `FDH2QHSX4_D_CP_SETUP_negedge_posedge, `FDH2QHSX4_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDH2QHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDH2QHSX4_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDH2QHSX4_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& D, `FDH2QHSX4_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D, posedge CD, `FDH2QHSX4_CD_CP_REM_posedge_posedge, Notifier);
 
`endif
   endspecify
`endif


endmodule // FDH2QHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:27 and Version :1.1 //
 
//  START 
// CELL FDH2QHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDH2QHSX8_CD_F_Q_F 0.1
`define FDH2QHSX8_CP_R_Q_R 0.1
`define FDH2QHSX8_CP_R_Q_F 0.1
`define FDH2QHSX8_D_CP_HOLD_posedge_posedge 0.1
`define FDH2QHSX8_D_CP_HOLD_negedge_posedge 0.1
`define FDH2QHSX8_D_CP_SETUP_posedge_posedge 0.1
`define FDH2QHSX8_D_CP_SETUP_negedge_posedge 0.1
`define FDH2QHSX8_CP_PWL 0.1
`define FDH2QHSX8_CP_PWH 0.1
`define FDH2QHSX8_CD_PWL 0.1
`define FDH2QHSX8_CD_CP_REC_posedge_posedge 0.1
`define FDH2QHSX8_CD_CP_REM_posedge_posedge 0.1

module FDH2QHSX8 (Q, D, CP, CD);

   output Q;
   input D;
   input CP;
   input CD;


   reg Notifier;


   U_FD_P_RN_NOTI u0 (IQ, D, CP, CD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(CD) (posedge CP => (Q +: D)) = (`FDH2QHSX8_CP_R_Q_R, `FDH2QHSX8_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FDH2QHSX8_CD_F_Q_F,`FDH2QHSX8_CD_F_Q_F);

	$setuphold(posedge CP &&& CD, posedge D, `FDH2QHSX8_D_CP_SETUP_posedge_posedge, `FDH2QHSX8_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge D, `FDH2QHSX8_D_CP_SETUP_negedge_posedge, `FDH2QHSX8_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDH2QHSX8_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDH2QHSX8_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDH2QHSX8_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& D, `FDH2QHSX8_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D, posedge CD, `FDH2QHSX8_CD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: D)) = (`FDH2QHSX8_CP_R_Q_R, `FDH2QHSX8_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FDH2QHSX8_CD_F_Q_F,`FDH2QHSX8_CD_F_Q_F);
 
        $setuphold(posedge CP &&& CD, posedge D, `FDH2QHSX8_D_CP_SETUP_posedge_posedge, `FDH2QHSX8_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge D, `FDH2QHSX8_D_CP_SETUP_negedge_posedge, `FDH2QHSX8_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDH2QHSX8_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDH2QHSX8_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDH2QHSX8_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& D, `FDH2QHSX8_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D, posedge CD, `FDH2QHSX8_CD_CP_REM_posedge_posedge, Notifier);
 
`endif
   endspecify
`endif


endmodule // FDH2QHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:27 and Version :1.1 //
 
//  START 
// CELL F_FD2QHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_FD2QHS_CD_F_Q_F 0.1
`define F_FD2QHS_CP_R_Q_R 0.1
`define F_FD2QHS_CP_R_Q_F 0.1
`define F_FD2QHS_D_CP_HOLD_posedge_posedge 0.1
`define F_FD2QHS_D_CP_HOLD_negedge_posedge 0.1
`define F_FD2QHS_D_CP_SETUP_posedge_posedge 0.1
`define F_FD2QHS_D_CP_SETUP_negedge_posedge 0.1
`define F_FD2QHS_CP_PWL 0.1
`define F_FD2QHS_CP_PWH 0.1
`define F_FD2QHS_CD_PWL 0.1
`define F_FD2QHS_CD_CP_REC_posedge_posedge 0.1
`define F_FD2QHS_CD_CP_REM_posedge_posedge 0.1

module F_FD2QHS (Q, D, CP, CD);

   output Q;
   input D;
   input CP;
   input CD;


   reg Notifier;


   U_FD_P_RN_NOTI u0 (IQ, D, CP, CD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(CD) (posedge CP => (Q +: D)) = (`F_FD2QHS_CP_R_Q_R, `F_FD2QHS_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`F_FD2QHS_CD_F_Q_F,`F_FD2QHS_CD_F_Q_F);

	$setuphold(posedge CP &&& CD, posedge D, `F_FD2QHS_D_CP_SETUP_posedge_posedge, `F_FD2QHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge D, `F_FD2QHS_D_CP_SETUP_negedge_posedge, `F_FD2QHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `F_FD2QHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `F_FD2QHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `F_FD2QHS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& D, `F_FD2QHS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D, posedge CD, `F_FD2QHS_CD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: D)) = (`F_FD2QHS_CP_R_Q_R, `F_FD2QHS_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`F_FD2QHS_CD_F_Q_F,`F_FD2QHS_CD_F_Q_F);
 
        $setuphold(posedge CP &&& CD, posedge D, `F_FD2QHS_D_CP_SETUP_posedge_posedge, `F_FD2QHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge D, `F_FD2QHS_D_CP_SETUP_negedge_posedge, `F_FD2QHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `F_FD2QHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `F_FD2QHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `F_FD2QHS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& D, `F_FD2QHS_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D, posedge CD, `F_FD2QHS_CD_CP_REM_posedge_posedge, Notifier);
 
`endif
   endspecify
`endif


endmodule // F_FD2QHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:27 and Version :1.1 //
 
//  START 
// CELL F_FD2QHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_FD2QHSP_CD_F_Q_F 0.1
`define F_FD2QHSP_CP_R_Q_R 0.1
`define F_FD2QHSP_CP_R_Q_F 0.1
`define F_FD2QHSP_D_CP_HOLD_posedge_posedge 0.1
`define F_FD2QHSP_D_CP_HOLD_negedge_posedge 0.1
`define F_FD2QHSP_D_CP_SETUP_posedge_posedge 0.1
`define F_FD2QHSP_D_CP_SETUP_negedge_posedge 0.1
`define F_FD2QHSP_CP_PWL 0.1
`define F_FD2QHSP_CP_PWH 0.1
`define F_FD2QHSP_CD_PWL 0.1
`define F_FD2QHSP_CD_CP_REC_posedge_posedge 0.1
`define F_FD2QHSP_CD_CP_REM_posedge_posedge 0.1

module F_FD2QHSP (Q, D, CP, CD);

   output Q;
   input D;
   input CP;
   input CD;


   reg Notifier;


   U_FD_P_RN_NOTI u0 (IQ, D, CP, CD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(CD) (posedge CP => (Q +: D)) = (`F_FD2QHSP_CP_R_Q_R, `F_FD2QHSP_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`F_FD2QHSP_CD_F_Q_F,`F_FD2QHSP_CD_F_Q_F);

	$setuphold(posedge CP &&& CD, posedge D, `F_FD2QHSP_D_CP_SETUP_posedge_posedge, `F_FD2QHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge D, `F_FD2QHSP_D_CP_SETUP_negedge_posedge, `F_FD2QHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `F_FD2QHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `F_FD2QHSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `F_FD2QHSP_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& D, `F_FD2QHSP_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D, posedge CD, `F_FD2QHSP_CD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: D)) = (`F_FD2QHSP_CP_R_Q_R, `F_FD2QHSP_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`F_FD2QHSP_CD_F_Q_F,`F_FD2QHSP_CD_F_Q_F);
 
        $setuphold(posedge CP &&& CD, posedge D, `F_FD2QHSP_D_CP_SETUP_posedge_posedge, `F_FD2QHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge D, `F_FD2QHSP_D_CP_SETUP_negedge_posedge, `F_FD2QHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `F_FD2QHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `F_FD2QHSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `F_FD2QHSP_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& D, `F_FD2QHSP_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D, posedge CD, `F_FD2QHSP_CD_CP_REM_posedge_posedge, Notifier);
 
`endif
   endspecify
`endif


endmodule // F_FD2QHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:27 and Version :1.1 //
 
//  START 
// CELL F_FD2QHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_FD2QHSX4_CD_F_Q_F 0.1
`define F_FD2QHSX4_CP_R_Q_R 0.1
`define F_FD2QHSX4_CP_R_Q_F 0.1
`define F_FD2QHSX4_D_CP_HOLD_posedge_posedge 0.1
`define F_FD2QHSX4_D_CP_HOLD_negedge_posedge 0.1
`define F_FD2QHSX4_D_CP_SETUP_posedge_posedge 0.1
`define F_FD2QHSX4_D_CP_SETUP_negedge_posedge 0.1
`define F_FD2QHSX4_CP_PWL 0.1
`define F_FD2QHSX4_CP_PWH 0.1
`define F_FD2QHSX4_CD_PWL 0.1
`define F_FD2QHSX4_CD_CP_REC_posedge_posedge 0.1
`define F_FD2QHSX4_CD_CP_REM_posedge_posedge 0.1

module F_FD2QHSX4 (Q, D, CP, CD);

   output Q;
   input D;
   input CP;
   input CD;


   reg Notifier;


   U_FD_P_RN_NOTI u0 (IQ, D, CP, CD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(CD) (posedge CP => (Q +: D)) = (`F_FD2QHSX4_CP_R_Q_R, `F_FD2QHSX4_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`F_FD2QHSX4_CD_F_Q_F,`F_FD2QHSX4_CD_F_Q_F);

	$setuphold(posedge CP &&& CD, posedge D, `F_FD2QHSX4_D_CP_SETUP_posedge_posedge, `F_FD2QHSX4_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge D, `F_FD2QHSX4_D_CP_SETUP_negedge_posedge, `F_FD2QHSX4_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `F_FD2QHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `F_FD2QHSX4_CP_PWH, 0, Notifier);
      $width(negedge CD, `F_FD2QHSX4_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& D, `F_FD2QHSX4_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D, posedge CD, `F_FD2QHSX4_CD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: D)) = (`F_FD2QHSX4_CP_R_Q_R, `F_FD2QHSX4_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`F_FD2QHSX4_CD_F_Q_F,`F_FD2QHSX4_CD_F_Q_F);
 
        $setuphold(posedge CP &&& CD, posedge D, `F_FD2QHSX4_D_CP_SETUP_posedge_posedge, `F_FD2QHSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge D, `F_FD2QHSX4_D_CP_SETUP_negedge_posedge, `F_FD2QHSX4_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `F_FD2QHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `F_FD2QHSX4_CP_PWH, 0, Notifier);
      $width(negedge CD, `F_FD2QHSX4_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& D, `F_FD2QHSX4_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D, posedge CD, `F_FD2QHSX4_CD_CP_REM_posedge_posedge, Notifier);
 
`endif
   endspecify
`endif


endmodule // F_FD2QHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:27 and Version :1.1 //
 
//  START 
// CELL FD2Q_SYNCHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD2Q_SYNCHS_NCD_R_Q_F 0.1
`define FD2Q_SYNCHS_CP_R_Q_R 0.1
`define FD2Q_SYNCHS_CP_R_Q_F 0.1
`define FD2Q_SYNCHS_D_CP_HOLD_posedge_posedge 0.1
`define FD2Q_SYNCHS_D_CP_HOLD_negedge_posedge 0.1
`define FD2Q_SYNCHS_D_CP_SETUP_posedge_posedge 0.1
`define FD2Q_SYNCHS_D_CP_SETUP_negedge_posedge 0.1
`define FD2Q_SYNCHS_CP_PWL 0.1
`define FD2Q_SYNCHS_CP_PWH 0.1
`define FD2Q_SYNCHS_NCD_PWH 0.1
`define FD2Q_SYNCHS_NCD_CP_REC_negedge_posedge 0.1
`define FD2Q_SYNCHS_NCD_CP_REM_negedge_posedge 0.1

module FD2Q_SYNCHS (Q, D, CP, NCD);

   output Q;
   input D;
   input CP;
   input NCD;


   reg Notifier;

   not u0 (CD, NCD);

   U_FD_P_RN_NOTI u1 (IQ, D, CP, CD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(CD) (posedge CP => (Q +: D)) = (`FD2Q_SYNCHS_CP_R_Q_R, `FD2Q_SYNCHS_CP_R_Q_F);
      (posedge NCD => (Q +: 1'b0)) = (`FD2Q_SYNCHS_NCD_R_Q_F,`FD2Q_SYNCHS_NCD_R_Q_F);

	$setuphold(posedge CP &&& CD, posedge D, `FD2Q_SYNCHS_D_CP_SETUP_posedge_posedge, `FD2Q_SYNCHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge D, `FD2Q_SYNCHS_D_CP_SETUP_negedge_posedge, `FD2Q_SYNCHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD2Q_SYNCHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2Q_SYNCHS_CP_PWH, 0, Notifier);
      $width(posedge NCD, `FD2Q_SYNCHS_NCD_PWH, 0, Notifier);

      $recovery(negedge NCD, posedge CP &&& D, `FD2Q_SYNCHS_NCD_CP_REC_negedge_posedge, Notifier);
      $hold(posedge CP &&& D, negedge NCD, `FD2Q_SYNCHS_NCD_CP_REM_negedge_posedge, Notifier);

`else

      (posedge CP => (Q +: D)) = (`FD2Q_SYNCHS_CP_R_Q_R, `FD2Q_SYNCHS_CP_R_Q_F);
      (posedge NCD => (Q +: 1'b0)) = (`FD2Q_SYNCHS_NCD_R_Q_F,`FD2Q_SYNCHS_NCD_R_Q_F);
 
        $setuphold(posedge CP &&& CD, posedge D, `FD2Q_SYNCHS_D_CP_SETUP_posedge_posedge, `FD2Q_SYNCHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge D, `FD2Q_SYNCHS_D_CP_SETUP_negedge_posedge, `FD2Q_SYNCHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD2Q_SYNCHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2Q_SYNCHS_CP_PWH, 0, Notifier);
      $width(posedge NCD, `FD2Q_SYNCHS_NCD_PWH, 0, Notifier);
 
      $recovery(negedge NCD, posedge CP &&& D, `FD2Q_SYNCHS_NCD_CP_REC_negedge_posedge, Notifier);
      $hold(posedge CP &&& D, negedge NCD, `FD2Q_SYNCHS_NCD_CP_REM_negedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FD2Q_SYNCHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:32 and Version :1.1 //
 
//  START 
// CELL FD2SHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD2SHS_CD_F_QN_R 0.1
`define FD2SHS_CP_R_QN_F 0.1
`define FD2SHS_CP_R_QN_R 0.1
`define FD2SHS_CD_F_Q_F 0.1
`define FD2SHS_CP_R_Q_R 0.1
`define FD2SHS_CP_R_Q_F 0.1
`define FD2SHS_CD_CP_REM_posedge_posedge 0.1
`define FD2SHS_CD_CP_REC_posedge_posedge 0.1
`define FD2SHS_CD_PWL 0.1
`define FD2SHS_CP_PWH 0.1
`define FD2SHS_CP_PWL 0.1
`define FD2SHS_D_CP_SETUP_posedge_posedge 0.1
`define FD2SHS_D_CP_SETUP_negedge_posedge 0.1
`define FD2SHS_D_CP_HOLD_posedge_posedge 0.1
`define FD2SHS_D_CP_HOLD_negedge_posedge 0.1
`define FD2SHS_TI_CP_SETUP_posedge_posedge 0.1
`define FD2SHS_TI_CP_SETUP_negedge_posedge 0.1
`define FD2SHS_TI_CP_HOLD_posedge_posedge 0.1
`define FD2SHS_TI_CP_HOLD_negedge_posedge 0.1
`define FD2SHS_TE_CP_SETUP_posedge_posedge 0.1
`define FD2SHS_TE_CP_SETUP_negedge_posedge 0.1
`define FD2SHS_TE_CP_HOLD_posedge_posedge 0.1
`define FD2SHS_TE_CP_HOLD_negedge_posedge 0.1

module FD2SHS (Q, QN, D, CP, CD, TI, TE);

   output Q;
   output QN;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);

   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && CD) (posedge CP => (Q +: D)) = (`FD2SHS_CP_R_Q_R, `FD2SHS_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`FD2SHS_CP_R_Q_R, `FD2SHS_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`FD2SHS_CP_R_Q_R, `FD2SHS_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`FD2SHS_CP_R_Q_R, `FD2SHS_CP_R_Q_F);
      if(!TE && CD) (posedge CP => (QN -: D)) = (`FD2SHS_CP_R_QN_R, `FD2SHS_CP_R_QN_F);
      if(TE && CD) (posedge CP => (QN -: TI)) = (`FD2SHS_CP_R_QN_R, `FD2SHS_CP_R_QN_F);
      if(!D && TI && CD) (posedge CP => (QN -: TE)) = (`FD2SHS_CP_R_QN_R, `FD2SHS_CP_R_QN_F);
      if(!TI && D && CD) (posedge CP => (QN +: TE)) = (`FD2SHS_CP_R_QN_R, `FD2SHS_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2SHS_CD_F_Q_F,`FD2SHS_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FD2SHS_CD_F_QN_R,`FD2SHS_CD_F_QN_R);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FD2SHS_TE_CP_SETUP_posedge_posedge, `FD2SHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FD2SHS_TE_CP_SETUP_negedge_posedge, `FD2SHS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `FD2SHS_TI_CP_SETUP_posedge_posedge, `FD2SHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `FD2SHS_TI_CP_SETUP_negedge_posedge, `FD2SHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `FD2SHS_D_CP_SETUP_posedge_posedge, `FD2SHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `FD2SHS_D_CP_SETUP_negedge_posedge, `FD2SHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD2SHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2SHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2SHS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FD2SHS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `FD2SHS_CD_CP_REM_posedge_posedge, Notifier);
`else 
       (posedge CP => (Q +: Mux21DTITE_)) = (`FD2SHS_CP_R_Q_R, `FD2SHS_CP_R_Q_F);
       (posedge CP => (QN -: Mux21DTITE_)) = (`FD2SHS_CP_R_QN_R, `FD2SHS_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2SHS_CD_F_Q_F,`FD2SHS_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FD2SHS_CD_F_QN_R,`FD2SHS_CD_F_QN_R);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FD2SHS_TE_CP_SETUP_posedge_posedge, `FD2SHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FD2SHS_TE_CP_SETUP_negedge_posedge, `FD2SHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `FD2SHS_TI_CP_SETUP_posedge_posedge,`FD2SHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `FD2SHS_TI_CP_SETUP_negedge_posedge,`FD2SHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `FD2SHS_D_CP_SETUP_posedge_posedge,`FD2SHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `FD2SHS_D_CP_SETUP_negedge_posedge,`FD2SHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD2SHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2SHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2SHS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FD2SHS_CD_CP_REC_posedge_posedge,Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `FD2SHS_CD_CP_REM_posedge_posedge, Notifier);


`endif

   endspecify
`endif


endmodule // FD2SHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:32 and Version :1.1 //
 
//  START 
// CELL FD2SHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD2SHSP_CD_F_QN_R 0.1
`define FD2SHSP_CP_R_QN_F 0.1
`define FD2SHSP_CP_R_QN_R 0.1
`define FD2SHSP_CD_F_Q_F 0.1
`define FD2SHSP_CP_R_Q_R 0.1
`define FD2SHSP_CP_R_Q_F 0.1
`define FD2SHSP_CD_CP_REM_posedge_posedge 0.1
`define FD2SHSP_CD_CP_REC_posedge_posedge 0.1
`define FD2SHSP_CD_PWL 0.1
`define FD2SHSP_CP_PWH 0.1
`define FD2SHSP_CP_PWL 0.1
`define FD2SHSP_D_CP_SETUP_posedge_posedge 0.1
`define FD2SHSP_D_CP_SETUP_negedge_posedge 0.1
`define FD2SHSP_D_CP_HOLD_posedge_posedge 0.1
`define FD2SHSP_D_CP_HOLD_negedge_posedge 0.1
`define FD2SHSP_TI_CP_SETUP_posedge_posedge 0.1
`define FD2SHSP_TI_CP_SETUP_negedge_posedge 0.1
`define FD2SHSP_TI_CP_HOLD_posedge_posedge 0.1
`define FD2SHSP_TI_CP_HOLD_negedge_posedge 0.1
`define FD2SHSP_TE_CP_SETUP_posedge_posedge 0.1
`define FD2SHSP_TE_CP_SETUP_negedge_posedge 0.1
`define FD2SHSP_TE_CP_HOLD_posedge_posedge 0.1
`define FD2SHSP_TE_CP_HOLD_negedge_posedge 0.1

module FD2SHSP (Q, QN, D, CP, CD, TI, TE);

   output Q;
   output QN;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);

   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && CD) (posedge CP => (Q +: D)) = (`FD2SHSP_CP_R_Q_R, `FD2SHSP_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`FD2SHSP_CP_R_Q_R, `FD2SHSP_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`FD2SHSP_CP_R_Q_R, `FD2SHSP_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`FD2SHSP_CP_R_Q_R, `FD2SHSP_CP_R_Q_F);
      if(!TE && CD) (posedge CP => (QN -: D)) = (`FD2SHSP_CP_R_QN_R, `FD2SHSP_CP_R_QN_F);
      if(TE && CD) (posedge CP => (QN -: TI)) = (`FD2SHSP_CP_R_QN_R, `FD2SHSP_CP_R_QN_F);
      if(!D && TI && CD) (posedge CP => (QN -: TE)) = (`FD2SHSP_CP_R_QN_R, `FD2SHSP_CP_R_QN_F);
      if(!TI && D && CD) (posedge CP => (QN +: TE)) = (`FD2SHSP_CP_R_QN_R, `FD2SHSP_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2SHSP_CD_F_Q_F,`FD2SHSP_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FD2SHSP_CD_F_QN_R,`FD2SHSP_CD_F_QN_R);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FD2SHSP_TE_CP_SETUP_posedge_posedge, `FD2SHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FD2SHSP_TE_CP_SETUP_negedge_posedge, `FD2SHSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `FD2SHSP_TI_CP_SETUP_posedge_posedge, `FD2SHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `FD2SHSP_TI_CP_SETUP_negedge_posedge, `FD2SHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `FD2SHSP_D_CP_SETUP_posedge_posedge, `FD2SHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `FD2SHSP_D_CP_SETUP_negedge_posedge, `FD2SHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD2SHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2SHSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2SHSP_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FD2SHSP_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `FD2SHSP_CD_CP_REM_posedge_posedge, Notifier);
`else 
       (posedge CP => (Q +: Mux21DTITE_)) = (`FD2SHSP_CP_R_Q_R, `FD2SHSP_CP_R_Q_F);
       (posedge CP => (QN -: Mux21DTITE_)) = (`FD2SHSP_CP_R_QN_R, `FD2SHSP_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2SHSP_CD_F_Q_F,`FD2SHSP_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FD2SHSP_CD_F_QN_R,`FD2SHSP_CD_F_QN_R);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FD2SHSP_TE_CP_SETUP_posedge_posedge, `FD2SHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FD2SHSP_TE_CP_SETUP_negedge_posedge, `FD2SHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `FD2SHSP_TI_CP_SETUP_posedge_posedge,`FD2SHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `FD2SHSP_TI_CP_SETUP_negedge_posedge,`FD2SHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `FD2SHSP_D_CP_SETUP_posedge_posedge,`FD2SHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `FD2SHSP_D_CP_SETUP_negedge_posedge,`FD2SHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD2SHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2SHSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2SHSP_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FD2SHSP_CD_CP_REC_posedge_posedge,Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `FD2SHSP_CD_CP_REM_posedge_posedge, Notifier);


`endif

   endspecify
`endif


endmodule // FD2SHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:32 and Version :1.1 //
 
//  START 
// CELL FDM2SHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDM2SHS_CD_F_QN_R 0.1
`define FDM2SHS_CP_R_QN_F 0.1
`define FDM2SHS_CP_R_QN_R 0.1
`define FDM2SHS_CD_F_Q_F 0.1
`define FDM2SHS_CP_R_Q_R 0.1
`define FDM2SHS_CP_R_Q_F 0.1
`define FDM2SHS_CD_CP_REM_posedge_posedge 0.1
`define FDM2SHS_CD_CP_REC_posedge_posedge 0.1
`define FDM2SHS_CD_PWL 0.1
`define FDM2SHS_CP_PWH 0.1
`define FDM2SHS_CP_PWL 0.1
`define FDM2SHS_D_CP_SETUP_posedge_posedge 0.1
`define FDM2SHS_D_CP_SETUP_negedge_posedge 0.1
`define FDM2SHS_D_CP_HOLD_posedge_posedge 0.1
`define FDM2SHS_D_CP_HOLD_negedge_posedge 0.1
`define FDM2SHS_TI_CP_SETUP_posedge_posedge 0.1
`define FDM2SHS_TI_CP_SETUP_negedge_posedge 0.1
`define FDM2SHS_TI_CP_HOLD_posedge_posedge 0.1
`define FDM2SHS_TI_CP_HOLD_negedge_posedge 0.1
`define FDM2SHS_TE_CP_SETUP_posedge_posedge 0.1
`define FDM2SHS_TE_CP_SETUP_negedge_posedge 0.1
`define FDM2SHS_TE_CP_HOLD_posedge_posedge 0.1
`define FDM2SHS_TE_CP_HOLD_negedge_posedge 0.1

module FDM2SHS (Q, QN, D, CP, CD, TI, TE);

   output Q;
   output QN;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);

   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && CD) (posedge CP => (Q +: D)) = (`FDM2SHS_CP_R_Q_R, `FDM2SHS_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`FDM2SHS_CP_R_Q_R, `FDM2SHS_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`FDM2SHS_CP_R_Q_R, `FDM2SHS_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`FDM2SHS_CP_R_Q_R, `FDM2SHS_CP_R_Q_F);
      if(!TE && CD) (posedge CP => (QN -: D)) = (`FDM2SHS_CP_R_QN_R, `FDM2SHS_CP_R_QN_F);
      if(TE && CD) (posedge CP => (QN -: TI)) = (`FDM2SHS_CP_R_QN_R, `FDM2SHS_CP_R_QN_F);
      if(!D && TI && CD) (posedge CP => (QN -: TE)) = (`FDM2SHS_CP_R_QN_R, `FDM2SHS_CP_R_QN_F);
      if(!TI && D && CD) (posedge CP => (QN +: TE)) = (`FDM2SHS_CP_R_QN_R, `FDM2SHS_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FDM2SHS_CD_F_Q_F,`FDM2SHS_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FDM2SHS_CD_F_QN_R,`FDM2SHS_CD_F_QN_R);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FDM2SHS_TE_CP_SETUP_posedge_posedge, `FDM2SHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FDM2SHS_TE_CP_SETUP_negedge_posedge, `FDM2SHS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `FDM2SHS_TI_CP_SETUP_posedge_posedge, `FDM2SHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `FDM2SHS_TI_CP_SETUP_negedge_posedge, `FDM2SHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `FDM2SHS_D_CP_SETUP_posedge_posedge, `FDM2SHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `FDM2SHS_D_CP_SETUP_negedge_posedge, `FDM2SHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDM2SHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDM2SHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDM2SHS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FDM2SHS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `FDM2SHS_CD_CP_REM_posedge_posedge, Notifier);
`else 
       (posedge CP => (Q +: Mux21DTITE_)) = (`FDM2SHS_CP_R_Q_R, `FDM2SHS_CP_R_Q_F);
       (posedge CP => (QN -: Mux21DTITE_)) = (`FDM2SHS_CP_R_QN_R, `FDM2SHS_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FDM2SHS_CD_F_Q_F,`FDM2SHS_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FDM2SHS_CD_F_QN_R,`FDM2SHS_CD_F_QN_R);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FDM2SHS_TE_CP_SETUP_posedge_posedge, `FDM2SHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FDM2SHS_TE_CP_SETUP_negedge_posedge, `FDM2SHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `FDM2SHS_TI_CP_SETUP_posedge_posedge,`FDM2SHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `FDM2SHS_TI_CP_SETUP_negedge_posedge,`FDM2SHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `FDM2SHS_D_CP_SETUP_posedge_posedge,`FDM2SHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `FDM2SHS_D_CP_SETUP_negedge_posedge,`FDM2SHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDM2SHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDM2SHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDM2SHS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FDM2SHS_CD_CP_REC_posedge_posedge,Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `FDM2SHS_CD_CP_REM_posedge_posedge, Notifier);


`endif

   endspecify
`endif


endmodule // FDM2SHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:32 and Version :1.1 //
 
//  START 
// CELL FDM2SHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDM2SHSP_CD_F_QN_R 0.1
`define FDM2SHSP_CP_R_QN_F 0.1
`define FDM2SHSP_CP_R_QN_R 0.1
`define FDM2SHSP_CD_F_Q_F 0.1
`define FDM2SHSP_CP_R_Q_R 0.1
`define FDM2SHSP_CP_R_Q_F 0.1
`define FDM2SHSP_CD_CP_REM_posedge_posedge 0.1
`define FDM2SHSP_CD_CP_REC_posedge_posedge 0.1
`define FDM2SHSP_CD_PWL 0.1
`define FDM2SHSP_CP_PWH 0.1
`define FDM2SHSP_CP_PWL 0.1
`define FDM2SHSP_D_CP_SETUP_posedge_posedge 0.1
`define FDM2SHSP_D_CP_SETUP_negedge_posedge 0.1
`define FDM2SHSP_D_CP_HOLD_posedge_posedge 0.1
`define FDM2SHSP_D_CP_HOLD_negedge_posedge 0.1
`define FDM2SHSP_TI_CP_SETUP_posedge_posedge 0.1
`define FDM2SHSP_TI_CP_SETUP_negedge_posedge 0.1
`define FDM2SHSP_TI_CP_HOLD_posedge_posedge 0.1
`define FDM2SHSP_TI_CP_HOLD_negedge_posedge 0.1
`define FDM2SHSP_TE_CP_SETUP_posedge_posedge 0.1
`define FDM2SHSP_TE_CP_SETUP_negedge_posedge 0.1
`define FDM2SHSP_TE_CP_HOLD_posedge_posedge 0.1
`define FDM2SHSP_TE_CP_HOLD_negedge_posedge 0.1

module FDM2SHSP (Q, QN, D, CP, CD, TI, TE);

   output Q;
   output QN;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);

   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && CD) (posedge CP => (Q +: D)) = (`FDM2SHSP_CP_R_Q_R, `FDM2SHSP_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`FDM2SHSP_CP_R_Q_R, `FDM2SHSP_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`FDM2SHSP_CP_R_Q_R, `FDM2SHSP_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`FDM2SHSP_CP_R_Q_R, `FDM2SHSP_CP_R_Q_F);
      if(!TE && CD) (posedge CP => (QN -: D)) = (`FDM2SHSP_CP_R_QN_R, `FDM2SHSP_CP_R_QN_F);
      if(TE && CD) (posedge CP => (QN -: TI)) = (`FDM2SHSP_CP_R_QN_R, `FDM2SHSP_CP_R_QN_F);
      if(!D && TI && CD) (posedge CP => (QN -: TE)) = (`FDM2SHSP_CP_R_QN_R, `FDM2SHSP_CP_R_QN_F);
      if(!TI && D && CD) (posedge CP => (QN +: TE)) = (`FDM2SHSP_CP_R_QN_R, `FDM2SHSP_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FDM2SHSP_CD_F_Q_F,`FDM2SHSP_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FDM2SHSP_CD_F_QN_R,`FDM2SHSP_CD_F_QN_R);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FDM2SHSP_TE_CP_SETUP_posedge_posedge, `FDM2SHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FDM2SHSP_TE_CP_SETUP_negedge_posedge, `FDM2SHSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `FDM2SHSP_TI_CP_SETUP_posedge_posedge, `FDM2SHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `FDM2SHSP_TI_CP_SETUP_negedge_posedge, `FDM2SHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `FDM2SHSP_D_CP_SETUP_posedge_posedge, `FDM2SHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `FDM2SHSP_D_CP_SETUP_negedge_posedge, `FDM2SHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDM2SHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDM2SHSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDM2SHSP_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FDM2SHSP_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `FDM2SHSP_CD_CP_REM_posedge_posedge, Notifier);
`else 
       (posedge CP => (Q +: Mux21DTITE_)) = (`FDM2SHSP_CP_R_Q_R, `FDM2SHSP_CP_R_Q_F);
       (posedge CP => (QN -: Mux21DTITE_)) = (`FDM2SHSP_CP_R_QN_R, `FDM2SHSP_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FDM2SHSP_CD_F_Q_F,`FDM2SHSP_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FDM2SHSP_CD_F_QN_R,`FDM2SHSP_CD_F_QN_R);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FDM2SHSP_TE_CP_SETUP_posedge_posedge, `FDM2SHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FDM2SHSP_TE_CP_SETUP_negedge_posedge, `FDM2SHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `FDM2SHSP_TI_CP_SETUP_posedge_posedge,`FDM2SHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `FDM2SHSP_TI_CP_SETUP_negedge_posedge,`FDM2SHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `FDM2SHSP_D_CP_SETUP_posedge_posedge,`FDM2SHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `FDM2SHSP_D_CP_SETUP_negedge_posedge,`FDM2SHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDM2SHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDM2SHSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDM2SHSP_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FDM2SHSP_CD_CP_REC_posedge_posedge,Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `FDM2SHSP_CD_CP_REM_posedge_posedge, Notifier);


`endif

   endspecify
`endif


endmodule // FDM2SHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:32 and Version :1.1 //
 
//  START 
// CELL FDH2SHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDH2SHSX4_CD_F_QN_R 0.1
`define FDH2SHSX4_CP_R_QN_F 0.1
`define FDH2SHSX4_CP_R_QN_R 0.1
`define FDH2SHSX4_CD_F_Q_F 0.1
`define FDH2SHSX4_CP_R_Q_R 0.1
`define FDH2SHSX4_CP_R_Q_F 0.1
`define FDH2SHSX4_CD_CP_REM_posedge_posedge 0.1
`define FDH2SHSX4_CD_CP_REC_posedge_posedge 0.1
`define FDH2SHSX4_CD_PWL 0.1
`define FDH2SHSX4_CP_PWH 0.1
`define FDH2SHSX4_CP_PWL 0.1
`define FDH2SHSX4_D_CP_SETUP_posedge_posedge 0.1
`define FDH2SHSX4_D_CP_SETUP_negedge_posedge 0.1
`define FDH2SHSX4_D_CP_HOLD_posedge_posedge 0.1
`define FDH2SHSX4_D_CP_HOLD_negedge_posedge 0.1
`define FDH2SHSX4_TI_CP_SETUP_posedge_posedge 0.1
`define FDH2SHSX4_TI_CP_SETUP_negedge_posedge 0.1
`define FDH2SHSX4_TI_CP_HOLD_posedge_posedge 0.1
`define FDH2SHSX4_TI_CP_HOLD_negedge_posedge 0.1
`define FDH2SHSX4_TE_CP_SETUP_posedge_posedge 0.1
`define FDH2SHSX4_TE_CP_SETUP_negedge_posedge 0.1
`define FDH2SHSX4_TE_CP_HOLD_posedge_posedge 0.1
`define FDH2SHSX4_TE_CP_HOLD_negedge_posedge 0.1

module FDH2SHSX4 (Q, QN, D, CP, CD, TI, TE);

   output Q;
   output QN;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);

   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && CD) (posedge CP => (Q +: D)) = (`FDH2SHSX4_CP_R_Q_R, `FDH2SHSX4_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`FDH2SHSX4_CP_R_Q_R, `FDH2SHSX4_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`FDH2SHSX4_CP_R_Q_R, `FDH2SHSX4_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`FDH2SHSX4_CP_R_Q_R, `FDH2SHSX4_CP_R_Q_F);
      if(!TE && CD) (posedge CP => (QN -: D)) = (`FDH2SHSX4_CP_R_QN_R, `FDH2SHSX4_CP_R_QN_F);
      if(TE && CD) (posedge CP => (QN -: TI)) = (`FDH2SHSX4_CP_R_QN_R, `FDH2SHSX4_CP_R_QN_F);
      if(!D && TI && CD) (posedge CP => (QN -: TE)) = (`FDH2SHSX4_CP_R_QN_R, `FDH2SHSX4_CP_R_QN_F);
      if(!TI && D && CD) (posedge CP => (QN +: TE)) = (`FDH2SHSX4_CP_R_QN_R, `FDH2SHSX4_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FDH2SHSX4_CD_F_Q_F,`FDH2SHSX4_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FDH2SHSX4_CD_F_QN_R,`FDH2SHSX4_CD_F_QN_R);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FDH2SHSX4_TE_CP_SETUP_posedge_posedge, `FDH2SHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FDH2SHSX4_TE_CP_SETUP_negedge_posedge, `FDH2SHSX4_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `FDH2SHSX4_TI_CP_SETUP_posedge_posedge, `FDH2SHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `FDH2SHSX4_TI_CP_SETUP_negedge_posedge, `FDH2SHSX4_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `FDH2SHSX4_D_CP_SETUP_posedge_posedge, `FDH2SHSX4_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `FDH2SHSX4_D_CP_SETUP_negedge_posedge, `FDH2SHSX4_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDH2SHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDH2SHSX4_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDH2SHSX4_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FDH2SHSX4_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `FDH2SHSX4_CD_CP_REM_posedge_posedge, Notifier);
`else 
       (posedge CP => (Q +: Mux21DTITE_)) = (`FDH2SHSX4_CP_R_Q_R, `FDH2SHSX4_CP_R_Q_F);
       (posedge CP => (QN -: Mux21DTITE_)) = (`FDH2SHSX4_CP_R_QN_R, `FDH2SHSX4_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FDH2SHSX4_CD_F_Q_F,`FDH2SHSX4_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FDH2SHSX4_CD_F_QN_R,`FDH2SHSX4_CD_F_QN_R);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FDH2SHSX4_TE_CP_SETUP_posedge_posedge, `FDH2SHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FDH2SHSX4_TE_CP_SETUP_negedge_posedge, `FDH2SHSX4_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `FDH2SHSX4_TI_CP_SETUP_posedge_posedge,`FDH2SHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `FDH2SHSX4_TI_CP_SETUP_negedge_posedge,`FDH2SHSX4_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `FDH2SHSX4_D_CP_SETUP_posedge_posedge,`FDH2SHSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `FDH2SHSX4_D_CP_SETUP_negedge_posedge,`FDH2SHSX4_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDH2SHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDH2SHSX4_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDH2SHSX4_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FDH2SHSX4_CD_CP_REC_posedge_posedge,Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `FDH2SHSX4_CD_CP_REM_posedge_posedge, Notifier);


`endif

   endspecify
`endif


endmodule // FDH2SHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:32 and Version :1.1 //
 
//  START 
// CELL FDH2SHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDH2SHSX8_CD_F_QN_R 0.1
`define FDH2SHSX8_CP_R_QN_F 0.1
`define FDH2SHSX8_CP_R_QN_R 0.1
`define FDH2SHSX8_CD_F_Q_F 0.1
`define FDH2SHSX8_CP_R_Q_R 0.1
`define FDH2SHSX8_CP_R_Q_F 0.1
`define FDH2SHSX8_CD_CP_REM_posedge_posedge 0.1
`define FDH2SHSX8_CD_CP_REC_posedge_posedge 0.1
`define FDH2SHSX8_CD_PWL 0.1
`define FDH2SHSX8_CP_PWH 0.1
`define FDH2SHSX8_CP_PWL 0.1
`define FDH2SHSX8_D_CP_SETUP_posedge_posedge 0.1
`define FDH2SHSX8_D_CP_SETUP_negedge_posedge 0.1
`define FDH2SHSX8_D_CP_HOLD_posedge_posedge 0.1
`define FDH2SHSX8_D_CP_HOLD_negedge_posedge 0.1
`define FDH2SHSX8_TI_CP_SETUP_posedge_posedge 0.1
`define FDH2SHSX8_TI_CP_SETUP_negedge_posedge 0.1
`define FDH2SHSX8_TI_CP_HOLD_posedge_posedge 0.1
`define FDH2SHSX8_TI_CP_HOLD_negedge_posedge 0.1
`define FDH2SHSX8_TE_CP_SETUP_posedge_posedge 0.1
`define FDH2SHSX8_TE_CP_SETUP_negedge_posedge 0.1
`define FDH2SHSX8_TE_CP_HOLD_posedge_posedge 0.1
`define FDH2SHSX8_TE_CP_HOLD_negedge_posedge 0.1

module FDH2SHSX8 (Q, QN, D, CP, CD, TI, TE);

   output Q;
   output QN;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);

   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && CD) (posedge CP => (Q +: D)) = (`FDH2SHSX8_CP_R_Q_R, `FDH2SHSX8_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`FDH2SHSX8_CP_R_Q_R, `FDH2SHSX8_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`FDH2SHSX8_CP_R_Q_R, `FDH2SHSX8_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`FDH2SHSX8_CP_R_Q_R, `FDH2SHSX8_CP_R_Q_F);
      if(!TE && CD) (posedge CP => (QN -: D)) = (`FDH2SHSX8_CP_R_QN_R, `FDH2SHSX8_CP_R_QN_F);
      if(TE && CD) (posedge CP => (QN -: TI)) = (`FDH2SHSX8_CP_R_QN_R, `FDH2SHSX8_CP_R_QN_F);
      if(!D && TI && CD) (posedge CP => (QN -: TE)) = (`FDH2SHSX8_CP_R_QN_R, `FDH2SHSX8_CP_R_QN_F);
      if(!TI && D && CD) (posedge CP => (QN +: TE)) = (`FDH2SHSX8_CP_R_QN_R, `FDH2SHSX8_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FDH2SHSX8_CD_F_Q_F,`FDH2SHSX8_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FDH2SHSX8_CD_F_QN_R,`FDH2SHSX8_CD_F_QN_R);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FDH2SHSX8_TE_CP_SETUP_posedge_posedge, `FDH2SHSX8_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FDH2SHSX8_TE_CP_SETUP_negedge_posedge, `FDH2SHSX8_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `FDH2SHSX8_TI_CP_SETUP_posedge_posedge, `FDH2SHSX8_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `FDH2SHSX8_TI_CP_SETUP_negedge_posedge, `FDH2SHSX8_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `FDH2SHSX8_D_CP_SETUP_posedge_posedge, `FDH2SHSX8_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `FDH2SHSX8_D_CP_SETUP_negedge_posedge, `FDH2SHSX8_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDH2SHSX8_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDH2SHSX8_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDH2SHSX8_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FDH2SHSX8_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `FDH2SHSX8_CD_CP_REM_posedge_posedge, Notifier);
`else 
       (posedge CP => (Q +: Mux21DTITE_)) = (`FDH2SHSX8_CP_R_Q_R, `FDH2SHSX8_CP_R_Q_F);
       (posedge CP => (QN -: Mux21DTITE_)) = (`FDH2SHSX8_CP_R_QN_R, `FDH2SHSX8_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FDH2SHSX8_CD_F_Q_F,`FDH2SHSX8_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FDH2SHSX8_CD_F_QN_R,`FDH2SHSX8_CD_F_QN_R);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FDH2SHSX8_TE_CP_SETUP_posedge_posedge, `FDH2SHSX8_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FDH2SHSX8_TE_CP_SETUP_negedge_posedge, `FDH2SHSX8_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `FDH2SHSX8_TI_CP_SETUP_posedge_posedge,`FDH2SHSX8_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `FDH2SHSX8_TI_CP_SETUP_negedge_posedge,`FDH2SHSX8_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `FDH2SHSX8_D_CP_SETUP_posedge_posedge,`FDH2SHSX8_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `FDH2SHSX8_D_CP_SETUP_negedge_posedge,`FDH2SHSX8_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDH2SHSX8_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDH2SHSX8_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDH2SHSX8_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FDH2SHSX8_CD_CP_REC_posedge_posedge,Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `FDH2SHSX8_CD_CP_REM_posedge_posedge, Notifier);


`endif

   endspecify
`endif


endmodule // FDH2SHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:32 and Version :1.1 //
 
//  START 
// CELL F_FD2SHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_FD2SHS_CD_F_QN_R 0.1
`define F_FD2SHS_CP_R_QN_F 0.1
`define F_FD2SHS_CP_R_QN_R 0.1
`define F_FD2SHS_CD_F_Q_F 0.1
`define F_FD2SHS_CP_R_Q_R 0.1
`define F_FD2SHS_CP_R_Q_F 0.1
`define F_FD2SHS_CD_CP_REM_posedge_posedge 0.1
`define F_FD2SHS_CD_CP_REC_posedge_posedge 0.1
`define F_FD2SHS_CD_PWL 0.1
`define F_FD2SHS_CP_PWH 0.1
`define F_FD2SHS_CP_PWL 0.1
`define F_FD2SHS_D_CP_SETUP_posedge_posedge 0.1
`define F_FD2SHS_D_CP_SETUP_negedge_posedge 0.1
`define F_FD2SHS_D_CP_HOLD_posedge_posedge 0.1
`define F_FD2SHS_D_CP_HOLD_negedge_posedge 0.1
`define F_FD2SHS_TI_CP_SETUP_posedge_posedge 0.1
`define F_FD2SHS_TI_CP_SETUP_negedge_posedge 0.1
`define F_FD2SHS_TI_CP_HOLD_posedge_posedge 0.1
`define F_FD2SHS_TI_CP_HOLD_negedge_posedge 0.1
`define F_FD2SHS_TE_CP_SETUP_posedge_posedge 0.1
`define F_FD2SHS_TE_CP_SETUP_negedge_posedge 0.1
`define F_FD2SHS_TE_CP_HOLD_posedge_posedge 0.1
`define F_FD2SHS_TE_CP_HOLD_negedge_posedge 0.1

module F_FD2SHS (Q, QN, D, CP, CD, TI, TE);

   output Q;
   output QN;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);

   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && CD) (posedge CP => (Q +: D)) = (`F_FD2SHS_CP_R_Q_R, `F_FD2SHS_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`F_FD2SHS_CP_R_Q_R, `F_FD2SHS_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`F_FD2SHS_CP_R_Q_R, `F_FD2SHS_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`F_FD2SHS_CP_R_Q_R, `F_FD2SHS_CP_R_Q_F);
      if(!TE && CD) (posedge CP => (QN -: D)) = (`F_FD2SHS_CP_R_QN_R, `F_FD2SHS_CP_R_QN_F);
      if(TE && CD) (posedge CP => (QN -: TI)) = (`F_FD2SHS_CP_R_QN_R, `F_FD2SHS_CP_R_QN_F);
      if(!D && TI && CD) (posedge CP => (QN -: TE)) = (`F_FD2SHS_CP_R_QN_R, `F_FD2SHS_CP_R_QN_F);
      if(!TI && D && CD) (posedge CP => (QN +: TE)) = (`F_FD2SHS_CP_R_QN_R, `F_FD2SHS_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`F_FD2SHS_CD_F_Q_F,`F_FD2SHS_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`F_FD2SHS_CD_F_QN_R,`F_FD2SHS_CD_F_QN_R);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `F_FD2SHS_TE_CP_SETUP_posedge_posedge, `F_FD2SHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `F_FD2SHS_TE_CP_SETUP_negedge_posedge, `F_FD2SHS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `F_FD2SHS_TI_CP_SETUP_posedge_posedge, `F_FD2SHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `F_FD2SHS_TI_CP_SETUP_negedge_posedge, `F_FD2SHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `F_FD2SHS_D_CP_SETUP_posedge_posedge, `F_FD2SHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `F_FD2SHS_D_CP_SETUP_negedge_posedge, `F_FD2SHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `F_FD2SHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `F_FD2SHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `F_FD2SHS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `F_FD2SHS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `F_FD2SHS_CD_CP_REM_posedge_posedge, Notifier);
`else 
       (posedge CP => (Q +: Mux21DTITE_)) = (`F_FD2SHS_CP_R_Q_R, `F_FD2SHS_CP_R_Q_F);
       (posedge CP => (QN -: Mux21DTITE_)) = (`F_FD2SHS_CP_R_QN_R, `F_FD2SHS_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`F_FD2SHS_CD_F_Q_F,`F_FD2SHS_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`F_FD2SHS_CD_F_QN_R,`F_FD2SHS_CD_F_QN_R);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `F_FD2SHS_TE_CP_SETUP_posedge_posedge, `F_FD2SHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `F_FD2SHS_TE_CP_SETUP_negedge_posedge, `F_FD2SHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `F_FD2SHS_TI_CP_SETUP_posedge_posedge,`F_FD2SHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `F_FD2SHS_TI_CP_SETUP_negedge_posedge,`F_FD2SHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `F_FD2SHS_D_CP_SETUP_posedge_posedge,`F_FD2SHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `F_FD2SHS_D_CP_SETUP_negedge_posedge,`F_FD2SHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `F_FD2SHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `F_FD2SHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `F_FD2SHS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `F_FD2SHS_CD_CP_REC_posedge_posedge,Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `F_FD2SHS_CD_CP_REM_posedge_posedge, Notifier);


`endif

   endspecify
`endif


endmodule // F_FD2SHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:32 and Version :1.1 //
 
//  START 
// CELL F_FD2SHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_FD2SHSP_CD_F_QN_R 0.1
`define F_FD2SHSP_CP_R_QN_F 0.1
`define F_FD2SHSP_CP_R_QN_R 0.1
`define F_FD2SHSP_CD_F_Q_F 0.1
`define F_FD2SHSP_CP_R_Q_R 0.1
`define F_FD2SHSP_CP_R_Q_F 0.1
`define F_FD2SHSP_CD_CP_REM_posedge_posedge 0.1
`define F_FD2SHSP_CD_CP_REC_posedge_posedge 0.1
`define F_FD2SHSP_CD_PWL 0.1
`define F_FD2SHSP_CP_PWH 0.1
`define F_FD2SHSP_CP_PWL 0.1
`define F_FD2SHSP_D_CP_SETUP_posedge_posedge 0.1
`define F_FD2SHSP_D_CP_SETUP_negedge_posedge 0.1
`define F_FD2SHSP_D_CP_HOLD_posedge_posedge 0.1
`define F_FD2SHSP_D_CP_HOLD_negedge_posedge 0.1
`define F_FD2SHSP_TI_CP_SETUP_posedge_posedge 0.1
`define F_FD2SHSP_TI_CP_SETUP_negedge_posedge 0.1
`define F_FD2SHSP_TI_CP_HOLD_posedge_posedge 0.1
`define F_FD2SHSP_TI_CP_HOLD_negedge_posedge 0.1
`define F_FD2SHSP_TE_CP_SETUP_posedge_posedge 0.1
`define F_FD2SHSP_TE_CP_SETUP_negedge_posedge 0.1
`define F_FD2SHSP_TE_CP_HOLD_posedge_posedge 0.1
`define F_FD2SHSP_TE_CP_HOLD_negedge_posedge 0.1

module F_FD2SHSP (Q, QN, D, CP, CD, TI, TE);

   output Q;
   output QN;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);

   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && CD) (posedge CP => (Q +: D)) = (`F_FD2SHSP_CP_R_Q_R, `F_FD2SHSP_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`F_FD2SHSP_CP_R_Q_R, `F_FD2SHSP_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`F_FD2SHSP_CP_R_Q_R, `F_FD2SHSP_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`F_FD2SHSP_CP_R_Q_R, `F_FD2SHSP_CP_R_Q_F);
      if(!TE && CD) (posedge CP => (QN -: D)) = (`F_FD2SHSP_CP_R_QN_R, `F_FD2SHSP_CP_R_QN_F);
      if(TE && CD) (posedge CP => (QN -: TI)) = (`F_FD2SHSP_CP_R_QN_R, `F_FD2SHSP_CP_R_QN_F);
      if(!D && TI && CD) (posedge CP => (QN -: TE)) = (`F_FD2SHSP_CP_R_QN_R, `F_FD2SHSP_CP_R_QN_F);
      if(!TI && D && CD) (posedge CP => (QN +: TE)) = (`F_FD2SHSP_CP_R_QN_R, `F_FD2SHSP_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`F_FD2SHSP_CD_F_Q_F,`F_FD2SHSP_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`F_FD2SHSP_CD_F_QN_R,`F_FD2SHSP_CD_F_QN_R);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `F_FD2SHSP_TE_CP_SETUP_posedge_posedge, `F_FD2SHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `F_FD2SHSP_TE_CP_SETUP_negedge_posedge, `F_FD2SHSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `F_FD2SHSP_TI_CP_SETUP_posedge_posedge, `F_FD2SHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `F_FD2SHSP_TI_CP_SETUP_negedge_posedge, `F_FD2SHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `F_FD2SHSP_D_CP_SETUP_posedge_posedge, `F_FD2SHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `F_FD2SHSP_D_CP_SETUP_negedge_posedge, `F_FD2SHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `F_FD2SHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `F_FD2SHSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `F_FD2SHSP_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `F_FD2SHSP_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `F_FD2SHSP_CD_CP_REM_posedge_posedge, Notifier);
`else 
       (posedge CP => (Q +: Mux21DTITE_)) = (`F_FD2SHSP_CP_R_Q_R, `F_FD2SHSP_CP_R_Q_F);
       (posedge CP => (QN -: Mux21DTITE_)) = (`F_FD2SHSP_CP_R_QN_R, `F_FD2SHSP_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`F_FD2SHSP_CD_F_Q_F,`F_FD2SHSP_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`F_FD2SHSP_CD_F_QN_R,`F_FD2SHSP_CD_F_QN_R);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `F_FD2SHSP_TE_CP_SETUP_posedge_posedge, `F_FD2SHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `F_FD2SHSP_TE_CP_SETUP_negedge_posedge, `F_FD2SHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `F_FD2SHSP_TI_CP_SETUP_posedge_posedge,`F_FD2SHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `F_FD2SHSP_TI_CP_SETUP_negedge_posedge,`F_FD2SHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `F_FD2SHSP_D_CP_SETUP_posedge_posedge,`F_FD2SHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `F_FD2SHSP_D_CP_SETUP_negedge_posedge,`F_FD2SHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `F_FD2SHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `F_FD2SHSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `F_FD2SHSP_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `F_FD2SHSP_CD_CP_REC_posedge_posedge,Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `F_FD2SHSP_CD_CP_REM_posedge_posedge, Notifier);


`endif

   endspecify
`endif


endmodule // F_FD2SHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:32 and Version :1.1 //
 
//  START 
// CELL FD2SQHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD2SQHS_CD_F_Q_F 0.1
`define FD2SQHS_CP_R_Q_R 0.1
`define FD2SQHS_CP_R_Q_F 0.1
`define FD2SQHS_TE_CP_HOLD_posedge_posedge 0.1
`define FD2SQHS_TE_CP_HOLD_negedge_posedge 0.1
`define FD2SQHS_TE_CP_SETUP_posedge_posedge 0.1
`define FD2SQHS_TE_CP_SETUP_negedge_posedge 0.1
`define FD2SQHS_TI_CP_HOLD_posedge_posedge 0.1
`define FD2SQHS_TI_CP_HOLD_negedge_posedge 0.1
`define FD2SQHS_TI_CP_SETUP_posedge_posedge 0.1
`define FD2SQHS_TI_CP_SETUP_negedge_posedge 0.1
`define FD2SQHS_D_CP_HOLD_posedge_posedge 0.1
`define FD2SQHS_D_CP_HOLD_negedge_posedge 0.1
`define FD2SQHS_D_CP_SETUP_posedge_posedge 0.1
`define FD2SQHS_D_CP_SETUP_negedge_posedge 0.1
`define FD2SQHS_CP_PWL 0.1
`define FD2SQHS_CP_PWH 0.1
`define FD2SQHS_CD_PWL 0.1
`define FD2SQHS_CD_CP_REC_posedge_posedge 0.1
`define FD2SQHS_CD_CP_REM_posedge_posedge 0.1

module FD2SQHS (Q, D, CP, CD, TI, TE);

   output Q;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);
 

   specify
`ifdef verifault 

      if(!TE && CD) (posedge CP => (Q +: D)) = (`FD2SQHS_CP_R_Q_R, `FD2SQHS_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`FD2SQHS_CP_R_Q_R, `FD2SQHS_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`FD2SQHS_CP_R_Q_R, `FD2SQHS_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`FD2SQHS_CP_R_Q_R, `FD2SQHS_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2SQHS_CD_F_Q_F,`FD2SQHS_CD_F_Q_F);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FD2SQHS_TE_CP_SETUP_posedge_posedge, `FD2SQHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FD2SQHS_TE_CP_SETUP_negedge_posedge, `FD2SQHS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `FD2SQHS_TI_CP_SETUP_posedge_posedge, `FD2SQHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `FD2SQHS_TI_CP_SETUP_negedge_posedge, `FD2SQHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `FD2SQHS_D_CP_SETUP_posedge_posedge, `FD2SQHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `FD2SQHS_D_CP_SETUP_negedge_posedge, `FD2SQHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD2SQHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2SQHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2SQHS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FD2SQHS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `FD2SQHS_CD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FD2SQHS_CP_R_Q_R, `FD2SQHS_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2SQHS_CD_F_Q_F,`FD2SQHS_CD_F_Q_F);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FD2SQHS_TE_CP_SETUP_posedge_posedge, `FD2SQHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FD2SQHS_TE_CP_SETUP_negedge_posedge, `FD2SQHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `FD2SQHS_TI_CP_SETUP_posedge_posedge, `FD2SQHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `FD2SQHS_TI_CP_SETUP_negedge_posedge, `FD2SQHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `FD2SQHS_D_CP_SETUP_posedge_posedge,`FD2SQHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `FD2SQHS_D_CP_SETUP_negedge_posedge,`FD2SQHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD2SQHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2SQHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2SQHS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FD2SQHS_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `FD2SQHS_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FD2SQHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:38 and Version :1.1 //
 
//  START 
// CELL FD2SQHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD2SQHSP_CD_F_Q_F 0.1
`define FD2SQHSP_CP_R_Q_R 0.1
`define FD2SQHSP_CP_R_Q_F 0.1
`define FD2SQHSP_TE_CP_HOLD_posedge_posedge 0.1
`define FD2SQHSP_TE_CP_HOLD_negedge_posedge 0.1
`define FD2SQHSP_TE_CP_SETUP_posedge_posedge 0.1
`define FD2SQHSP_TE_CP_SETUP_negedge_posedge 0.1
`define FD2SQHSP_TI_CP_HOLD_posedge_posedge 0.1
`define FD2SQHSP_TI_CP_HOLD_negedge_posedge 0.1
`define FD2SQHSP_TI_CP_SETUP_posedge_posedge 0.1
`define FD2SQHSP_TI_CP_SETUP_negedge_posedge 0.1
`define FD2SQHSP_D_CP_HOLD_posedge_posedge 0.1
`define FD2SQHSP_D_CP_HOLD_negedge_posedge 0.1
`define FD2SQHSP_D_CP_SETUP_posedge_posedge 0.1
`define FD2SQHSP_D_CP_SETUP_negedge_posedge 0.1
`define FD2SQHSP_CP_PWL 0.1
`define FD2SQHSP_CP_PWH 0.1
`define FD2SQHSP_CD_PWL 0.1
`define FD2SQHSP_CD_CP_REC_posedge_posedge 0.1
`define FD2SQHSP_CD_CP_REM_posedge_posedge 0.1

module FD2SQHSP (Q, D, CP, CD, TI, TE);

   output Q;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);
 

   specify
`ifdef verifault 

      if(!TE && CD) (posedge CP => (Q +: D)) = (`FD2SQHSP_CP_R_Q_R, `FD2SQHSP_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`FD2SQHSP_CP_R_Q_R, `FD2SQHSP_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`FD2SQHSP_CP_R_Q_R, `FD2SQHSP_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`FD2SQHSP_CP_R_Q_R, `FD2SQHSP_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2SQHSP_CD_F_Q_F,`FD2SQHSP_CD_F_Q_F);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FD2SQHSP_TE_CP_SETUP_posedge_posedge, `FD2SQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FD2SQHSP_TE_CP_SETUP_negedge_posedge, `FD2SQHSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `FD2SQHSP_TI_CP_SETUP_posedge_posedge, `FD2SQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `FD2SQHSP_TI_CP_SETUP_negedge_posedge, `FD2SQHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `FD2SQHSP_D_CP_SETUP_posedge_posedge, `FD2SQHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `FD2SQHSP_D_CP_SETUP_negedge_posedge, `FD2SQHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD2SQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2SQHSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2SQHSP_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FD2SQHSP_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `FD2SQHSP_CD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FD2SQHSP_CP_R_Q_R, `FD2SQHSP_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2SQHSP_CD_F_Q_F,`FD2SQHSP_CD_F_Q_F);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FD2SQHSP_TE_CP_SETUP_posedge_posedge, `FD2SQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FD2SQHSP_TE_CP_SETUP_negedge_posedge, `FD2SQHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `FD2SQHSP_TI_CP_SETUP_posedge_posedge, `FD2SQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `FD2SQHSP_TI_CP_SETUP_negedge_posedge, `FD2SQHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `FD2SQHSP_D_CP_SETUP_posedge_posedge,`FD2SQHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `FD2SQHSP_D_CP_SETUP_negedge_posedge,`FD2SQHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD2SQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2SQHSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2SQHSP_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FD2SQHSP_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `FD2SQHSP_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FD2SQHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:38 and Version :1.1 //
 
//  START 
// CELL FD2SQHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD2SQHSX4_CD_F_Q_F 0.1
`define FD2SQHSX4_CP_R_Q_R 0.1
`define FD2SQHSX4_CP_R_Q_F 0.1
`define FD2SQHSX4_TE_CP_HOLD_posedge_posedge 0.1
`define FD2SQHSX4_TE_CP_HOLD_negedge_posedge 0.1
`define FD2SQHSX4_TE_CP_SETUP_posedge_posedge 0.1
`define FD2SQHSX4_TE_CP_SETUP_negedge_posedge 0.1
`define FD2SQHSX4_TI_CP_HOLD_posedge_posedge 0.1
`define FD2SQHSX4_TI_CP_HOLD_negedge_posedge 0.1
`define FD2SQHSX4_TI_CP_SETUP_posedge_posedge 0.1
`define FD2SQHSX4_TI_CP_SETUP_negedge_posedge 0.1
`define FD2SQHSX4_D_CP_HOLD_posedge_posedge 0.1
`define FD2SQHSX4_D_CP_HOLD_negedge_posedge 0.1
`define FD2SQHSX4_D_CP_SETUP_posedge_posedge 0.1
`define FD2SQHSX4_D_CP_SETUP_negedge_posedge 0.1
`define FD2SQHSX4_CP_PWL 0.1
`define FD2SQHSX4_CP_PWH 0.1
`define FD2SQHSX4_CD_PWL 0.1
`define FD2SQHSX4_CD_CP_REC_posedge_posedge 0.1
`define FD2SQHSX4_CD_CP_REM_posedge_posedge 0.1

module FD2SQHSX4 (Q, D, CP, CD, TI, TE);

   output Q;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);
 

   specify
`ifdef verifault 

      if(!TE && CD) (posedge CP => (Q +: D)) = (`FD2SQHSX4_CP_R_Q_R, `FD2SQHSX4_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`FD2SQHSX4_CP_R_Q_R, `FD2SQHSX4_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`FD2SQHSX4_CP_R_Q_R, `FD2SQHSX4_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`FD2SQHSX4_CP_R_Q_R, `FD2SQHSX4_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2SQHSX4_CD_F_Q_F,`FD2SQHSX4_CD_F_Q_F);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FD2SQHSX4_TE_CP_SETUP_posedge_posedge, `FD2SQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FD2SQHSX4_TE_CP_SETUP_negedge_posedge, `FD2SQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `FD2SQHSX4_TI_CP_SETUP_posedge_posedge, `FD2SQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `FD2SQHSX4_TI_CP_SETUP_negedge_posedge, `FD2SQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `FD2SQHSX4_D_CP_SETUP_posedge_posedge, `FD2SQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `FD2SQHSX4_D_CP_SETUP_negedge_posedge, `FD2SQHSX4_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD2SQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2SQHSX4_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2SQHSX4_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FD2SQHSX4_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `FD2SQHSX4_CD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FD2SQHSX4_CP_R_Q_R, `FD2SQHSX4_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2SQHSX4_CD_F_Q_F,`FD2SQHSX4_CD_F_Q_F);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FD2SQHSX4_TE_CP_SETUP_posedge_posedge, `FD2SQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FD2SQHSX4_TE_CP_SETUP_negedge_posedge, `FD2SQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `FD2SQHSX4_TI_CP_SETUP_posedge_posedge, `FD2SQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `FD2SQHSX4_TI_CP_SETUP_negedge_posedge, `FD2SQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `FD2SQHSX4_D_CP_SETUP_posedge_posedge,`FD2SQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `FD2SQHSX4_D_CP_SETUP_negedge_posedge,`FD2SQHSX4_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD2SQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2SQHSX4_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2SQHSX4_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FD2SQHSX4_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `FD2SQHSX4_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FD2SQHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:38 and Version :1.1 //
 
//  START 
// CELL FDM2SQHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDM2SQHS_CD_F_Q_F 0.1
`define FDM2SQHS_CP_R_Q_R 0.1
`define FDM2SQHS_CP_R_Q_F 0.1
`define FDM2SQHS_TE_CP_HOLD_posedge_posedge 0.1
`define FDM2SQHS_TE_CP_HOLD_negedge_posedge 0.1
`define FDM2SQHS_TE_CP_SETUP_posedge_posedge 0.1
`define FDM2SQHS_TE_CP_SETUP_negedge_posedge 0.1
`define FDM2SQHS_TI_CP_HOLD_posedge_posedge 0.1
`define FDM2SQHS_TI_CP_HOLD_negedge_posedge 0.1
`define FDM2SQHS_TI_CP_SETUP_posedge_posedge 0.1
`define FDM2SQHS_TI_CP_SETUP_negedge_posedge 0.1
`define FDM2SQHS_D_CP_HOLD_posedge_posedge 0.1
`define FDM2SQHS_D_CP_HOLD_negedge_posedge 0.1
`define FDM2SQHS_D_CP_SETUP_posedge_posedge 0.1
`define FDM2SQHS_D_CP_SETUP_negedge_posedge 0.1
`define FDM2SQHS_CP_PWL 0.1
`define FDM2SQHS_CP_PWH 0.1
`define FDM2SQHS_CD_PWL 0.1
`define FDM2SQHS_CD_CP_REC_posedge_posedge 0.1
`define FDM2SQHS_CD_CP_REM_posedge_posedge 0.1

module FDM2SQHS (Q, D, CP, CD, TI, TE);

   output Q;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);
 

   specify
`ifdef verifault 

      if(!TE && CD) (posedge CP => (Q +: D)) = (`FDM2SQHS_CP_R_Q_R, `FDM2SQHS_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`FDM2SQHS_CP_R_Q_R, `FDM2SQHS_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`FDM2SQHS_CP_R_Q_R, `FDM2SQHS_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`FDM2SQHS_CP_R_Q_R, `FDM2SQHS_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FDM2SQHS_CD_F_Q_F,`FDM2SQHS_CD_F_Q_F);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FDM2SQHS_TE_CP_SETUP_posedge_posedge, `FDM2SQHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FDM2SQHS_TE_CP_SETUP_negedge_posedge, `FDM2SQHS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `FDM2SQHS_TI_CP_SETUP_posedge_posedge, `FDM2SQHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `FDM2SQHS_TI_CP_SETUP_negedge_posedge, `FDM2SQHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `FDM2SQHS_D_CP_SETUP_posedge_posedge, `FDM2SQHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `FDM2SQHS_D_CP_SETUP_negedge_posedge, `FDM2SQHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDM2SQHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDM2SQHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDM2SQHS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FDM2SQHS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `FDM2SQHS_CD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FDM2SQHS_CP_R_Q_R, `FDM2SQHS_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FDM2SQHS_CD_F_Q_F,`FDM2SQHS_CD_F_Q_F);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FDM2SQHS_TE_CP_SETUP_posedge_posedge, `FDM2SQHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FDM2SQHS_TE_CP_SETUP_negedge_posedge, `FDM2SQHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `FDM2SQHS_TI_CP_SETUP_posedge_posedge, `FDM2SQHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `FDM2SQHS_TI_CP_SETUP_negedge_posedge, `FDM2SQHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `FDM2SQHS_D_CP_SETUP_posedge_posedge,`FDM2SQHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `FDM2SQHS_D_CP_SETUP_negedge_posedge,`FDM2SQHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDM2SQHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDM2SQHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDM2SQHS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FDM2SQHS_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `FDM2SQHS_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FDM2SQHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:38 and Version :1.1 //
 
//  START 
// CELL FDM2SQHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDM2SQHSP_CD_F_Q_F 0.1
`define FDM2SQHSP_CP_R_Q_R 0.1
`define FDM2SQHSP_CP_R_Q_F 0.1
`define FDM2SQHSP_TE_CP_HOLD_posedge_posedge 0.1
`define FDM2SQHSP_TE_CP_HOLD_negedge_posedge 0.1
`define FDM2SQHSP_TE_CP_SETUP_posedge_posedge 0.1
`define FDM2SQHSP_TE_CP_SETUP_negedge_posedge 0.1
`define FDM2SQHSP_TI_CP_HOLD_posedge_posedge 0.1
`define FDM2SQHSP_TI_CP_HOLD_negedge_posedge 0.1
`define FDM2SQHSP_TI_CP_SETUP_posedge_posedge 0.1
`define FDM2SQHSP_TI_CP_SETUP_negedge_posedge 0.1
`define FDM2SQHSP_D_CP_HOLD_posedge_posedge 0.1
`define FDM2SQHSP_D_CP_HOLD_negedge_posedge 0.1
`define FDM2SQHSP_D_CP_SETUP_posedge_posedge 0.1
`define FDM2SQHSP_D_CP_SETUP_negedge_posedge 0.1
`define FDM2SQHSP_CP_PWL 0.1
`define FDM2SQHSP_CP_PWH 0.1
`define FDM2SQHSP_CD_PWL 0.1
`define FDM2SQHSP_CD_CP_REC_posedge_posedge 0.1
`define FDM2SQHSP_CD_CP_REM_posedge_posedge 0.1

module FDM2SQHSP (Q, D, CP, CD, TI, TE);

   output Q;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);
 

   specify
`ifdef verifault 

      if(!TE && CD) (posedge CP => (Q +: D)) = (`FDM2SQHSP_CP_R_Q_R, `FDM2SQHSP_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`FDM2SQHSP_CP_R_Q_R, `FDM2SQHSP_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`FDM2SQHSP_CP_R_Q_R, `FDM2SQHSP_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`FDM2SQHSP_CP_R_Q_R, `FDM2SQHSP_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FDM2SQHSP_CD_F_Q_F,`FDM2SQHSP_CD_F_Q_F);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FDM2SQHSP_TE_CP_SETUP_posedge_posedge, `FDM2SQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FDM2SQHSP_TE_CP_SETUP_negedge_posedge, `FDM2SQHSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `FDM2SQHSP_TI_CP_SETUP_posedge_posedge, `FDM2SQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `FDM2SQHSP_TI_CP_SETUP_negedge_posedge, `FDM2SQHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `FDM2SQHSP_D_CP_SETUP_posedge_posedge, `FDM2SQHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `FDM2SQHSP_D_CP_SETUP_negedge_posedge, `FDM2SQHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDM2SQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDM2SQHSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDM2SQHSP_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FDM2SQHSP_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `FDM2SQHSP_CD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FDM2SQHSP_CP_R_Q_R, `FDM2SQHSP_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FDM2SQHSP_CD_F_Q_F,`FDM2SQHSP_CD_F_Q_F);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FDM2SQHSP_TE_CP_SETUP_posedge_posedge, `FDM2SQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FDM2SQHSP_TE_CP_SETUP_negedge_posedge, `FDM2SQHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `FDM2SQHSP_TI_CP_SETUP_posedge_posedge, `FDM2SQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `FDM2SQHSP_TI_CP_SETUP_negedge_posedge, `FDM2SQHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `FDM2SQHSP_D_CP_SETUP_posedge_posedge,`FDM2SQHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `FDM2SQHSP_D_CP_SETUP_negedge_posedge,`FDM2SQHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDM2SQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDM2SQHSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDM2SQHSP_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FDM2SQHSP_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `FDM2SQHSP_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FDM2SQHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:38 and Version :1.1 //
 
//  START 
// CELL FDH2SQHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDH2SQHSX4_CD_F_Q_F 0.1
`define FDH2SQHSX4_CP_R_Q_R 0.1
`define FDH2SQHSX4_CP_R_Q_F 0.1
`define FDH2SQHSX4_TE_CP_HOLD_posedge_posedge 0.1
`define FDH2SQHSX4_TE_CP_HOLD_negedge_posedge 0.1
`define FDH2SQHSX4_TE_CP_SETUP_posedge_posedge 0.1
`define FDH2SQHSX4_TE_CP_SETUP_negedge_posedge 0.1
`define FDH2SQHSX4_TI_CP_HOLD_posedge_posedge 0.1
`define FDH2SQHSX4_TI_CP_HOLD_negedge_posedge 0.1
`define FDH2SQHSX4_TI_CP_SETUP_posedge_posedge 0.1
`define FDH2SQHSX4_TI_CP_SETUP_negedge_posedge 0.1
`define FDH2SQHSX4_D_CP_HOLD_posedge_posedge 0.1
`define FDH2SQHSX4_D_CP_HOLD_negedge_posedge 0.1
`define FDH2SQHSX4_D_CP_SETUP_posedge_posedge 0.1
`define FDH2SQHSX4_D_CP_SETUP_negedge_posedge 0.1
`define FDH2SQHSX4_CP_PWL 0.1
`define FDH2SQHSX4_CP_PWH 0.1
`define FDH2SQHSX4_CD_PWL 0.1
`define FDH2SQHSX4_CD_CP_REC_posedge_posedge 0.1
`define FDH2SQHSX4_CD_CP_REM_posedge_posedge 0.1

module FDH2SQHSX4 (Q, D, CP, CD, TI, TE);

   output Q;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);
 

   specify
`ifdef verifault 

      if(!TE && CD) (posedge CP => (Q +: D)) = (`FDH2SQHSX4_CP_R_Q_R, `FDH2SQHSX4_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`FDH2SQHSX4_CP_R_Q_R, `FDH2SQHSX4_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`FDH2SQHSX4_CP_R_Q_R, `FDH2SQHSX4_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`FDH2SQHSX4_CP_R_Q_R, `FDH2SQHSX4_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FDH2SQHSX4_CD_F_Q_F,`FDH2SQHSX4_CD_F_Q_F);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FDH2SQHSX4_TE_CP_SETUP_posedge_posedge, `FDH2SQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FDH2SQHSX4_TE_CP_SETUP_negedge_posedge, `FDH2SQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `FDH2SQHSX4_TI_CP_SETUP_posedge_posedge, `FDH2SQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `FDH2SQHSX4_TI_CP_SETUP_negedge_posedge, `FDH2SQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `FDH2SQHSX4_D_CP_SETUP_posedge_posedge, `FDH2SQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `FDH2SQHSX4_D_CP_SETUP_negedge_posedge, `FDH2SQHSX4_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDH2SQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDH2SQHSX4_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDH2SQHSX4_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FDH2SQHSX4_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `FDH2SQHSX4_CD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FDH2SQHSX4_CP_R_Q_R, `FDH2SQHSX4_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FDH2SQHSX4_CD_F_Q_F,`FDH2SQHSX4_CD_F_Q_F);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FDH2SQHSX4_TE_CP_SETUP_posedge_posedge, `FDH2SQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FDH2SQHSX4_TE_CP_SETUP_negedge_posedge, `FDH2SQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `FDH2SQHSX4_TI_CP_SETUP_posedge_posedge, `FDH2SQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `FDH2SQHSX4_TI_CP_SETUP_negedge_posedge, `FDH2SQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `FDH2SQHSX4_D_CP_SETUP_posedge_posedge,`FDH2SQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `FDH2SQHSX4_D_CP_SETUP_negedge_posedge,`FDH2SQHSX4_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDH2SQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDH2SQHSX4_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDH2SQHSX4_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FDH2SQHSX4_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `FDH2SQHSX4_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FDH2SQHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:38 and Version :1.1 //
 
//  START 
// CELL FDH2SQHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDH2SQHSX8_CD_F_Q_F 0.1
`define FDH2SQHSX8_CP_R_Q_R 0.1
`define FDH2SQHSX8_CP_R_Q_F 0.1
`define FDH2SQHSX8_TE_CP_HOLD_posedge_posedge 0.1
`define FDH2SQHSX8_TE_CP_HOLD_negedge_posedge 0.1
`define FDH2SQHSX8_TE_CP_SETUP_posedge_posedge 0.1
`define FDH2SQHSX8_TE_CP_SETUP_negedge_posedge 0.1
`define FDH2SQHSX8_TI_CP_HOLD_posedge_posedge 0.1
`define FDH2SQHSX8_TI_CP_HOLD_negedge_posedge 0.1
`define FDH2SQHSX8_TI_CP_SETUP_posedge_posedge 0.1
`define FDH2SQHSX8_TI_CP_SETUP_negedge_posedge 0.1
`define FDH2SQHSX8_D_CP_HOLD_posedge_posedge 0.1
`define FDH2SQHSX8_D_CP_HOLD_negedge_posedge 0.1
`define FDH2SQHSX8_D_CP_SETUP_posedge_posedge 0.1
`define FDH2SQHSX8_D_CP_SETUP_negedge_posedge 0.1
`define FDH2SQHSX8_CP_PWL 0.1
`define FDH2SQHSX8_CP_PWH 0.1
`define FDH2SQHSX8_CD_PWL 0.1
`define FDH2SQHSX8_CD_CP_REC_posedge_posedge 0.1
`define FDH2SQHSX8_CD_CP_REM_posedge_posedge 0.1

module FDH2SQHSX8 (Q, D, CP, CD, TI, TE);

   output Q;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);
 

   specify
`ifdef verifault 

      if(!TE && CD) (posedge CP => (Q +: D)) = (`FDH2SQHSX8_CP_R_Q_R, `FDH2SQHSX8_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`FDH2SQHSX8_CP_R_Q_R, `FDH2SQHSX8_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`FDH2SQHSX8_CP_R_Q_R, `FDH2SQHSX8_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`FDH2SQHSX8_CP_R_Q_R, `FDH2SQHSX8_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FDH2SQHSX8_CD_F_Q_F,`FDH2SQHSX8_CD_F_Q_F);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FDH2SQHSX8_TE_CP_SETUP_posedge_posedge, `FDH2SQHSX8_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FDH2SQHSX8_TE_CP_SETUP_negedge_posedge, `FDH2SQHSX8_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `FDH2SQHSX8_TI_CP_SETUP_posedge_posedge, `FDH2SQHSX8_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `FDH2SQHSX8_TI_CP_SETUP_negedge_posedge, `FDH2SQHSX8_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `FDH2SQHSX8_D_CP_SETUP_posedge_posedge, `FDH2SQHSX8_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `FDH2SQHSX8_D_CP_SETUP_negedge_posedge, `FDH2SQHSX8_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDH2SQHSX8_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDH2SQHSX8_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDH2SQHSX8_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FDH2SQHSX8_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `FDH2SQHSX8_CD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FDH2SQHSX8_CP_R_Q_R, `FDH2SQHSX8_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FDH2SQHSX8_CD_F_Q_F,`FDH2SQHSX8_CD_F_Q_F);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FDH2SQHSX8_TE_CP_SETUP_posedge_posedge, `FDH2SQHSX8_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FDH2SQHSX8_TE_CP_SETUP_negedge_posedge, `FDH2SQHSX8_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `FDH2SQHSX8_TI_CP_SETUP_posedge_posedge, `FDH2SQHSX8_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `FDH2SQHSX8_TI_CP_SETUP_negedge_posedge, `FDH2SQHSX8_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `FDH2SQHSX8_D_CP_SETUP_posedge_posedge,`FDH2SQHSX8_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `FDH2SQHSX8_D_CP_SETUP_negedge_posedge,`FDH2SQHSX8_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDH2SQHSX8_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDH2SQHSX8_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDH2SQHSX8_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FDH2SQHSX8_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `FDH2SQHSX8_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FDH2SQHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:38 and Version :1.1 //
 
//  START 
// CELL F_FD2SQHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_FD2SQHS_CD_F_Q_F 0.1
`define F_FD2SQHS_CP_R_Q_R 0.1
`define F_FD2SQHS_CP_R_Q_F 0.1
`define F_FD2SQHS_TE_CP_HOLD_posedge_posedge 0.1
`define F_FD2SQHS_TE_CP_HOLD_negedge_posedge 0.1
`define F_FD2SQHS_TE_CP_SETUP_posedge_posedge 0.1
`define F_FD2SQHS_TE_CP_SETUP_negedge_posedge 0.1
`define F_FD2SQHS_TI_CP_HOLD_posedge_posedge 0.1
`define F_FD2SQHS_TI_CP_HOLD_negedge_posedge 0.1
`define F_FD2SQHS_TI_CP_SETUP_posedge_posedge 0.1
`define F_FD2SQHS_TI_CP_SETUP_negedge_posedge 0.1
`define F_FD2SQHS_D_CP_HOLD_posedge_posedge 0.1
`define F_FD2SQHS_D_CP_HOLD_negedge_posedge 0.1
`define F_FD2SQHS_D_CP_SETUP_posedge_posedge 0.1
`define F_FD2SQHS_D_CP_SETUP_negedge_posedge 0.1
`define F_FD2SQHS_CP_PWL 0.1
`define F_FD2SQHS_CP_PWH 0.1
`define F_FD2SQHS_CD_PWL 0.1
`define F_FD2SQHS_CD_CP_REC_posedge_posedge 0.1
`define F_FD2SQHS_CD_CP_REM_posedge_posedge 0.1

module F_FD2SQHS (Q, D, CP, CD, TI, TE);

   output Q;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);
 

   specify
`ifdef verifault 

      if(!TE && CD) (posedge CP => (Q +: D)) = (`F_FD2SQHS_CP_R_Q_R, `F_FD2SQHS_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`F_FD2SQHS_CP_R_Q_R, `F_FD2SQHS_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`F_FD2SQHS_CP_R_Q_R, `F_FD2SQHS_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`F_FD2SQHS_CP_R_Q_R, `F_FD2SQHS_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`F_FD2SQHS_CD_F_Q_F,`F_FD2SQHS_CD_F_Q_F);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `F_FD2SQHS_TE_CP_SETUP_posedge_posedge, `F_FD2SQHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `F_FD2SQHS_TE_CP_SETUP_negedge_posedge, `F_FD2SQHS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `F_FD2SQHS_TI_CP_SETUP_posedge_posedge, `F_FD2SQHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `F_FD2SQHS_TI_CP_SETUP_negedge_posedge, `F_FD2SQHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `F_FD2SQHS_D_CP_SETUP_posedge_posedge, `F_FD2SQHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `F_FD2SQHS_D_CP_SETUP_negedge_posedge, `F_FD2SQHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `F_FD2SQHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `F_FD2SQHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `F_FD2SQHS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `F_FD2SQHS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `F_FD2SQHS_CD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`F_FD2SQHS_CP_R_Q_R, `F_FD2SQHS_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`F_FD2SQHS_CD_F_Q_F,`F_FD2SQHS_CD_F_Q_F);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `F_FD2SQHS_TE_CP_SETUP_posedge_posedge, `F_FD2SQHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `F_FD2SQHS_TE_CP_SETUP_negedge_posedge, `F_FD2SQHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `F_FD2SQHS_TI_CP_SETUP_posedge_posedge, `F_FD2SQHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `F_FD2SQHS_TI_CP_SETUP_negedge_posedge, `F_FD2SQHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `F_FD2SQHS_D_CP_SETUP_posedge_posedge,`F_FD2SQHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `F_FD2SQHS_D_CP_SETUP_negedge_posedge,`F_FD2SQHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `F_FD2SQHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `F_FD2SQHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `F_FD2SQHS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `F_FD2SQHS_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `F_FD2SQHS_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // F_FD2SQHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:38 and Version :1.1 //
 
//  START 
// CELL F_FD2SQHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_FD2SQHSP_CD_F_Q_F 0.1
`define F_FD2SQHSP_CP_R_Q_R 0.1
`define F_FD2SQHSP_CP_R_Q_F 0.1
`define F_FD2SQHSP_TE_CP_HOLD_posedge_posedge 0.1
`define F_FD2SQHSP_TE_CP_HOLD_negedge_posedge 0.1
`define F_FD2SQHSP_TE_CP_SETUP_posedge_posedge 0.1
`define F_FD2SQHSP_TE_CP_SETUP_negedge_posedge 0.1
`define F_FD2SQHSP_TI_CP_HOLD_posedge_posedge 0.1
`define F_FD2SQHSP_TI_CP_HOLD_negedge_posedge 0.1
`define F_FD2SQHSP_TI_CP_SETUP_posedge_posedge 0.1
`define F_FD2SQHSP_TI_CP_SETUP_negedge_posedge 0.1
`define F_FD2SQHSP_D_CP_HOLD_posedge_posedge 0.1
`define F_FD2SQHSP_D_CP_HOLD_negedge_posedge 0.1
`define F_FD2SQHSP_D_CP_SETUP_posedge_posedge 0.1
`define F_FD2SQHSP_D_CP_SETUP_negedge_posedge 0.1
`define F_FD2SQHSP_CP_PWL 0.1
`define F_FD2SQHSP_CP_PWH 0.1
`define F_FD2SQHSP_CD_PWL 0.1
`define F_FD2SQHSP_CD_CP_REC_posedge_posedge 0.1
`define F_FD2SQHSP_CD_CP_REM_posedge_posedge 0.1

module F_FD2SQHSP (Q, D, CP, CD, TI, TE);

   output Q;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);
 

   specify
`ifdef verifault 

      if(!TE && CD) (posedge CP => (Q +: D)) = (`F_FD2SQHSP_CP_R_Q_R, `F_FD2SQHSP_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`F_FD2SQHSP_CP_R_Q_R, `F_FD2SQHSP_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`F_FD2SQHSP_CP_R_Q_R, `F_FD2SQHSP_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`F_FD2SQHSP_CP_R_Q_R, `F_FD2SQHSP_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`F_FD2SQHSP_CD_F_Q_F,`F_FD2SQHSP_CD_F_Q_F);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `F_FD2SQHSP_TE_CP_SETUP_posedge_posedge, `F_FD2SQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `F_FD2SQHSP_TE_CP_SETUP_negedge_posedge, `F_FD2SQHSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `F_FD2SQHSP_TI_CP_SETUP_posedge_posedge, `F_FD2SQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `F_FD2SQHSP_TI_CP_SETUP_negedge_posedge, `F_FD2SQHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `F_FD2SQHSP_D_CP_SETUP_posedge_posedge, `F_FD2SQHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `F_FD2SQHSP_D_CP_SETUP_negedge_posedge, `F_FD2SQHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `F_FD2SQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `F_FD2SQHSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `F_FD2SQHSP_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `F_FD2SQHSP_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `F_FD2SQHSP_CD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`F_FD2SQHSP_CP_R_Q_R, `F_FD2SQHSP_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`F_FD2SQHSP_CD_F_Q_F,`F_FD2SQHSP_CD_F_Q_F);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `F_FD2SQHSP_TE_CP_SETUP_posedge_posedge, `F_FD2SQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `F_FD2SQHSP_TE_CP_SETUP_negedge_posedge, `F_FD2SQHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `F_FD2SQHSP_TI_CP_SETUP_posedge_posedge, `F_FD2SQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `F_FD2SQHSP_TI_CP_SETUP_negedge_posedge, `F_FD2SQHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `F_FD2SQHSP_D_CP_SETUP_posedge_posedge,`F_FD2SQHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `F_FD2SQHSP_D_CP_SETUP_negedge_posedge,`F_FD2SQHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `F_FD2SQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `F_FD2SQHSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `F_FD2SQHSP_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `F_FD2SQHSP_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `F_FD2SQHSP_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // F_FD2SQHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:38 and Version :1.1 //
 
//  START 
// CELL F_FD2SQHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_FD2SQHSX4_CD_F_Q_F 0.1
`define F_FD2SQHSX4_CP_R_Q_R 0.1
`define F_FD2SQHSX4_CP_R_Q_F 0.1
`define F_FD2SQHSX4_TE_CP_HOLD_posedge_posedge 0.1
`define F_FD2SQHSX4_TE_CP_HOLD_negedge_posedge 0.1
`define F_FD2SQHSX4_TE_CP_SETUP_posedge_posedge 0.1
`define F_FD2SQHSX4_TE_CP_SETUP_negedge_posedge 0.1
`define F_FD2SQHSX4_TI_CP_HOLD_posedge_posedge 0.1
`define F_FD2SQHSX4_TI_CP_HOLD_negedge_posedge 0.1
`define F_FD2SQHSX4_TI_CP_SETUP_posedge_posedge 0.1
`define F_FD2SQHSX4_TI_CP_SETUP_negedge_posedge 0.1
`define F_FD2SQHSX4_D_CP_HOLD_posedge_posedge 0.1
`define F_FD2SQHSX4_D_CP_HOLD_negedge_posedge 0.1
`define F_FD2SQHSX4_D_CP_SETUP_posedge_posedge 0.1
`define F_FD2SQHSX4_D_CP_SETUP_negedge_posedge 0.1
`define F_FD2SQHSX4_CP_PWL 0.1
`define F_FD2SQHSX4_CP_PWH 0.1
`define F_FD2SQHSX4_CD_PWL 0.1
`define F_FD2SQHSX4_CD_CP_REC_posedge_posedge 0.1
`define F_FD2SQHSX4_CD_CP_REM_posedge_posedge 0.1

module F_FD2SQHSX4 (Q, D, CP, CD, TI, TE);

   output Q;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);
 

   specify
`ifdef verifault 

      if(!TE && CD) (posedge CP => (Q +: D)) = (`F_FD2SQHSX4_CP_R_Q_R, `F_FD2SQHSX4_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`F_FD2SQHSX4_CP_R_Q_R, `F_FD2SQHSX4_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`F_FD2SQHSX4_CP_R_Q_R, `F_FD2SQHSX4_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`F_FD2SQHSX4_CP_R_Q_R, `F_FD2SQHSX4_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`F_FD2SQHSX4_CD_F_Q_F,`F_FD2SQHSX4_CD_F_Q_F);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `F_FD2SQHSX4_TE_CP_SETUP_posedge_posedge, `F_FD2SQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `F_FD2SQHSX4_TE_CP_SETUP_negedge_posedge, `F_FD2SQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `F_FD2SQHSX4_TI_CP_SETUP_posedge_posedge, `F_FD2SQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `F_FD2SQHSX4_TI_CP_SETUP_negedge_posedge, `F_FD2SQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `F_FD2SQHSX4_D_CP_SETUP_posedge_posedge, `F_FD2SQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `F_FD2SQHSX4_D_CP_SETUP_negedge_posedge, `F_FD2SQHSX4_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `F_FD2SQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `F_FD2SQHSX4_CP_PWH, 0, Notifier);
      $width(negedge CD, `F_FD2SQHSX4_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `F_FD2SQHSX4_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `F_FD2SQHSX4_CD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`F_FD2SQHSX4_CP_R_Q_R, `F_FD2SQHSX4_CP_R_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`F_FD2SQHSX4_CD_F_Q_F,`F_FD2SQHSX4_CD_F_Q_F);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `F_FD2SQHSX4_TE_CP_SETUP_posedge_posedge, `F_FD2SQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `F_FD2SQHSX4_TE_CP_SETUP_negedge_posedge, `F_FD2SQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `F_FD2SQHSX4_TI_CP_SETUP_posedge_posedge, `F_FD2SQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `F_FD2SQHSX4_TI_CP_SETUP_negedge_posedge, `F_FD2SQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `F_FD2SQHSX4_D_CP_SETUP_posedge_posedge,`F_FD2SQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `F_FD2SQHSX4_D_CP_SETUP_negedge_posedge,`F_FD2SQHSX4_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `F_FD2SQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `F_FD2SQHSX4_CP_PWH, 0, Notifier);
      $width(negedge CD, `F_FD2SQHSX4_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `F_FD2SQHSX4_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `F_FD2SQHSX4_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // F_FD2SQHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:38 and Version :1.1 //
 
//  START 
// CELL FD2THS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD2THS_CD_F_SO_F 0.1
`define FD2THS_CP_R_SO_R 0.1
`define FD2THS_CP_R_SO_F 0.1
`define FD2THS_CD_F_QN_R 0.1
`define FD2THS_CP_R_QN_F 0.1
`define FD2THS_CP_R_QN_R 0.1
`define FD2THS_CD_F_Q_F 0.1
`define FD2THS_CP_R_Q_R 0.1
`define FD2THS_CP_R_Q_F 0.1
`define FD2THS_CD_CP_REM_posedge_posedge 0.1
`define FD2THS_CD_CP_REC_posedge_posedge 0.1
`define FD2THS_CD_PWL 0.1
`define FD2THS_CP_PWH 0.1
`define FD2THS_CP_PWL 0.1
`define FD2THS_D_CP_SETUP_posedge_posedge 0.1
`define FD2THS_D_CP_SETUP_negedge_posedge 0.1
`define FD2THS_D_CP_HOLD_posedge_posedge 0.1
`define FD2THS_D_CP_HOLD_negedge_posedge 0.1
`define FD2THS_TI_CP_SETUP_posedge_posedge 0.1
`define FD2THS_TI_CP_SETUP_negedge_posedge 0.1
`define FD2THS_TI_CP_HOLD_posedge_posedge 0.1
`define FD2THS_TI_CP_HOLD_negedge_posedge 0.1
`define FD2THS_TE_CP_SETUP_posedge_posedge 0.1
`define FD2THS_TE_CP_SETUP_negedge_posedge 0.1
`define FD2THS_TE_CP_HOLD_posedge_posedge 0.1
`define FD2THS_TE_CP_HOLD_negedge_posedge 0.1

module FD2THS (Q, QN, SO, D, CP, CD, TI, TE);

   output Q;
   output QN;
   output SO;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);
   buf  u3 (SO, IQ);
   not  u4 (QN, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   and  (AndCDTEX_, CD, TEX);
   and  (AndCDTE_, CD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && CD) (posedge CP => (Q +: D)) = (`FD2THS_CP_R_Q_R, `FD2THS_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`FD2THS_CP_R_Q_R, `FD2THS_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`FD2THS_CP_R_Q_R, `FD2THS_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`FD2THS_CP_R_Q_R, `FD2THS_CP_R_Q_F);
      if(!TE && CD) (posedge CP => (QN -: D)) = (`FD2THS_CP_R_QN_R, `FD2THS_CP_R_QN_F);
      if(TE && CD) (posedge CP => (QN -: TI)) = (`FD2THS_CP_R_QN_R, `FD2THS_CP_R_QN_F);
      if(!D && TI && CD) (posedge CP => (QN -: TE)) = (`FD2THS_CP_R_QN_R, `FD2THS_CP_R_QN_F);
      if(!TI && D && CD) (posedge CP => (QN +: TE)) = (`FD2THS_CP_R_QN_R, `FD2THS_CP_R_QN_F);
      if(!TE && CD) (posedge CP => (SO +: D)) = (`FD2THS_CP_R_SO_R, `FD2THS_CP_R_SO_F);
      if(TE && CD) (posedge CP => (SO +: TI)) = (`FD2THS_CP_R_SO_R, `FD2THS_CP_R_SO_F);
      if(!D && TI && CD) (posedge CP => (SO +: TE)) = (`FD2THS_CP_R_SO_R, `FD2THS_CP_R_SO_F);
      if(!TI && D && CD) (posedge CP => (SO -: TE)) = (`FD2THS_CP_R_SO_R, `FD2THS_CP_R_SO_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2THS_CD_F_Q_F,`FD2THS_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FD2THS_CD_F_QN_R,`FD2THS_CD_F_QN_R);
      (negedge CD => (SO +: 1'b0)) = (`FD2THS_CD_F_SO_F,`FD2THS_CD_F_SO_F);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FD2THS_TE_CP_SETUP_posedge_posedge, `FD2THS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FD2THS_TE_CP_SETUP_negedge_posedge, `FD2THS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `FD2THS_TI_CP_SETUP_posedge_posedge, `FD2THS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `FD2THS_TI_CP_SETUP_negedge_posedge, `FD2THS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `FD2THS_D_CP_SETUP_posedge_posedge, `FD2THS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `FD2THS_D_CP_SETUP_negedge_posedge, `FD2THS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD2THS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2THS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2THS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FD2THS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `FD2THS_CD_CP_REM_posedge_posedge, Notifier);

`else

      (posedge CP => (Q +: Mux21DTITE_)) = (`FD2THS_CP_R_Q_R, `FD2THS_CP_R_Q_F);
      (posedge CP => (QN -: Mux21DTITE_)) = (`FD2THS_CP_R_QN_R, `FD2THS_CP_R_QN_F);
      (posedge CP => (SO +: Mux21DTITE_)) = (`FD2THS_CP_R_SO_R, `FD2THS_CP_R_SO_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2THS_CD_F_Q_F,`FD2THS_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FD2THS_CD_F_QN_R,`FD2THS_CD_F_QN_R);
      (negedge CD => (SO +: 1'b0)) = (`FD2THS_CD_F_SO_F,`FD2THS_CD_F_SO_F);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FD2THS_TE_CP_SETUP_posedge_posedge, `FD2THS_TE_CP_HOLD_posedge_posedge,Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FD2THS_TE_CP_SETUP_negedge_posedge, `FD2THS_TE_CP_HOLD_negedge_posedge,Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `FD2THS_TI_CP_SETUP_posedge_posedge, `FD2THS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `FD2THS_TI_CP_SETUP_negedge_posedge, `FD2THS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `FD2THS_D_CP_SETUP_posedge_posedge, `FD2THS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `FD2THS_D_CP_SETUP_negedge_posedge, `FD2THS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD2THS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2THS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2THS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FD2THS_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `FD2THS_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FD2THS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:45 and Version :1.1 //
 
//  START 
// CELL FD2THSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD2THSP_CD_F_SO_F 0.1
`define FD2THSP_CP_R_SO_R 0.1
`define FD2THSP_CP_R_SO_F 0.1
`define FD2THSP_CD_F_QN_R 0.1
`define FD2THSP_CP_R_QN_F 0.1
`define FD2THSP_CP_R_QN_R 0.1
`define FD2THSP_CD_F_Q_F 0.1
`define FD2THSP_CP_R_Q_R 0.1
`define FD2THSP_CP_R_Q_F 0.1
`define FD2THSP_CD_CP_REM_posedge_posedge 0.1
`define FD2THSP_CD_CP_REC_posedge_posedge 0.1
`define FD2THSP_CD_PWL 0.1
`define FD2THSP_CP_PWH 0.1
`define FD2THSP_CP_PWL 0.1
`define FD2THSP_D_CP_SETUP_posedge_posedge 0.1
`define FD2THSP_D_CP_SETUP_negedge_posedge 0.1
`define FD2THSP_D_CP_HOLD_posedge_posedge 0.1
`define FD2THSP_D_CP_HOLD_negedge_posedge 0.1
`define FD2THSP_TI_CP_SETUP_posedge_posedge 0.1
`define FD2THSP_TI_CP_SETUP_negedge_posedge 0.1
`define FD2THSP_TI_CP_HOLD_posedge_posedge 0.1
`define FD2THSP_TI_CP_HOLD_negedge_posedge 0.1
`define FD2THSP_TE_CP_SETUP_posedge_posedge 0.1
`define FD2THSP_TE_CP_SETUP_negedge_posedge 0.1
`define FD2THSP_TE_CP_HOLD_posedge_posedge 0.1
`define FD2THSP_TE_CP_HOLD_negedge_posedge 0.1

module FD2THSP (Q, QN, SO, D, CP, CD, TI, TE);

   output Q;
   output QN;
   output SO;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);
   buf  u3 (SO, IQ);
   not  u4 (QN, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   and  (AndCDTEX_, CD, TEX);
   and  (AndCDTE_, CD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && CD) (posedge CP => (Q +: D)) = (`FD2THSP_CP_R_Q_R, `FD2THSP_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`FD2THSP_CP_R_Q_R, `FD2THSP_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`FD2THSP_CP_R_Q_R, `FD2THSP_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`FD2THSP_CP_R_Q_R, `FD2THSP_CP_R_Q_F);
      if(!TE && CD) (posedge CP => (QN -: D)) = (`FD2THSP_CP_R_QN_R, `FD2THSP_CP_R_QN_F);
      if(TE && CD) (posedge CP => (QN -: TI)) = (`FD2THSP_CP_R_QN_R, `FD2THSP_CP_R_QN_F);
      if(!D && TI && CD) (posedge CP => (QN -: TE)) = (`FD2THSP_CP_R_QN_R, `FD2THSP_CP_R_QN_F);
      if(!TI && D && CD) (posedge CP => (QN +: TE)) = (`FD2THSP_CP_R_QN_R, `FD2THSP_CP_R_QN_F);
      if(!TE && CD) (posedge CP => (SO +: D)) = (`FD2THSP_CP_R_SO_R, `FD2THSP_CP_R_SO_F);
      if(TE && CD) (posedge CP => (SO +: TI)) = (`FD2THSP_CP_R_SO_R, `FD2THSP_CP_R_SO_F);
      if(!D && TI && CD) (posedge CP => (SO +: TE)) = (`FD2THSP_CP_R_SO_R, `FD2THSP_CP_R_SO_F);
      if(!TI && D && CD) (posedge CP => (SO -: TE)) = (`FD2THSP_CP_R_SO_R, `FD2THSP_CP_R_SO_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2THSP_CD_F_Q_F,`FD2THSP_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FD2THSP_CD_F_QN_R,`FD2THSP_CD_F_QN_R);
      (negedge CD => (SO +: 1'b0)) = (`FD2THSP_CD_F_SO_F,`FD2THSP_CD_F_SO_F);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FD2THSP_TE_CP_SETUP_posedge_posedge, `FD2THSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FD2THSP_TE_CP_SETUP_negedge_posedge, `FD2THSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `FD2THSP_TI_CP_SETUP_posedge_posedge, `FD2THSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `FD2THSP_TI_CP_SETUP_negedge_posedge, `FD2THSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `FD2THSP_D_CP_SETUP_posedge_posedge, `FD2THSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `FD2THSP_D_CP_SETUP_negedge_posedge, `FD2THSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD2THSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2THSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2THSP_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FD2THSP_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `FD2THSP_CD_CP_REM_posedge_posedge, Notifier);

`else

      (posedge CP => (Q +: Mux21DTITE_)) = (`FD2THSP_CP_R_Q_R, `FD2THSP_CP_R_Q_F);
      (posedge CP => (QN -: Mux21DTITE_)) = (`FD2THSP_CP_R_QN_R, `FD2THSP_CP_R_QN_F);
      (posedge CP => (SO +: Mux21DTITE_)) = (`FD2THSP_CP_R_SO_R, `FD2THSP_CP_R_SO_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2THSP_CD_F_Q_F,`FD2THSP_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FD2THSP_CD_F_QN_R,`FD2THSP_CD_F_QN_R);
      (negedge CD => (SO +: 1'b0)) = (`FD2THSP_CD_F_SO_F,`FD2THSP_CD_F_SO_F);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FD2THSP_TE_CP_SETUP_posedge_posedge, `FD2THSP_TE_CP_HOLD_posedge_posedge,Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FD2THSP_TE_CP_SETUP_negedge_posedge, `FD2THSP_TE_CP_HOLD_negedge_posedge,Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `FD2THSP_TI_CP_SETUP_posedge_posedge, `FD2THSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `FD2THSP_TI_CP_SETUP_negedge_posedge, `FD2THSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `FD2THSP_D_CP_SETUP_posedge_posedge, `FD2THSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `FD2THSP_D_CP_SETUP_negedge_posedge, `FD2THSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD2THSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2THSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2THSP_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FD2THSP_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `FD2THSP_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FD2THSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:45 and Version :1.1 //
 
//  START 
// CELL FD2TQHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD2TQHS_CD_F_SO_F 0.1
`define FD2TQHS_CP_R_SO_R 0.1
`define FD2TQHS_CP_R_SO_F 0.1
`define FD2TQHS_CD_F_Q_F 0.1
`define FD2TQHS_CP_R_Q_R 0.1
`define FD2TQHS_CP_R_Q_F 0.1
`define FD2TQHS_CD_CP_REM_posedge_posedge 0.1
`define FD2TQHS_CD_CP_REC_posedge_posedge 0.1
`define FD2TQHS_CD_PWL 0.1
`define FD2TQHS_CP_PWH 0.1
`define FD2TQHS_CP_PWL 0.1
`define FD2TQHS_D_CP_SETUP_posedge_posedge 0.1
`define FD2TQHS_D_CP_SETUP_negedge_posedge 0.1
`define FD2TQHS_D_CP_HOLD_posedge_posedge 0.1
`define FD2TQHS_D_CP_HOLD_negedge_posedge 0.1
`define FD2TQHS_TI_CP_SETUP_posedge_posedge 0.1
`define FD2TQHS_TI_CP_SETUP_negedge_posedge 0.1
`define FD2TQHS_TI_CP_HOLD_posedge_posedge 0.1
`define FD2TQHS_TI_CP_HOLD_negedge_posedge 0.1
`define FD2TQHS_TE_CP_SETUP_posedge_posedge 0.1
`define FD2TQHS_TE_CP_SETUP_negedge_posedge 0.1
`define FD2TQHS_TE_CP_HOLD_posedge_posedge 0.1
`define FD2TQHS_TE_CP_HOLD_negedge_posedge 0.1

module FD2TQHS (Q, SO, D, CP, CD, TI, TE);

   output Q;
   output SO;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);
   buf  u3 (SO, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   and  (AndCDTEX_, CD, TEX);
   and  (AndCDTE_, CD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && CD) (posedge CP => (Q +: D)) = (`FD2TQHS_CP_R_Q_R, `FD2TQHS_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`FD2TQHS_CP_R_Q_R, `FD2TQHS_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`FD2TQHS_CP_R_Q_R, `FD2TQHS_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`FD2TQHS_CP_R_Q_R, `FD2TQHS_CP_R_Q_F);
      if(!TE && CD) (posedge CP => (SO +: D)) = (`FD2TQHS_CP_R_SO_R, `FD2TQHS_CP_R_SO_F);
      if(TE && CD) (posedge CP => (SO +: TI)) = (`FD2TQHS_CP_R_SO_R, `FD2TQHS_CP_R_SO_F);
      if(!D && TI && CD) (posedge CP => (SO +: TE)) = (`FD2TQHS_CP_R_SO_R, `FD2TQHS_CP_R_SO_F);
      if(!TI && D && CD) (posedge CP => (SO -: TE)) = (`FD2TQHS_CP_R_SO_R, `FD2TQHS_CP_R_SO_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2TQHS_CD_F_Q_F,`FD2TQHS_CD_F_Q_F);
      (negedge CD => (SO +: 1'b0)) = (`FD2TQHS_CD_F_SO_F,`FD2TQHS_CD_F_SO_F);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FD2TQHS_TE_CP_SETUP_posedge_posedge, `FD2TQHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FD2TQHS_TE_CP_SETUP_negedge_posedge, `FD2TQHS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `FD2TQHS_TI_CP_SETUP_posedge_posedge, `FD2TQHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `FD2TQHS_TI_CP_SETUP_negedge_posedge, `FD2TQHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `FD2TQHS_D_CP_SETUP_posedge_posedge, `FD2TQHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `FD2TQHS_D_CP_SETUP_negedge_posedge, `FD2TQHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD2TQHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2TQHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2TQHS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FD2TQHS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `FD2TQHS_CD_CP_REM_posedge_posedge, Notifier);

`else
  (posedge CP => (Q +: Mux21DTITE_)) = (`FD2TQHS_CP_R_Q_R, `FD2TQHS_CP_R_Q_F);
      (posedge CP => (SO +: Mux21DTITE_)) = (`FD2TQHS_CP_R_SO_R, `FD2TQHS_CP_R_SO_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2TQHS_CD_F_Q_F,`FD2TQHS_CD_F_Q_F);
      (negedge CD => (SO +: 1'b0)) = (`FD2TQHS_CD_F_SO_F,`FD2TQHS_CD_F_SO_F);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FD2TQHS_TE_CP_SETUP_posedge_posedge, `FD2TQHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FD2TQHS_TE_CP_SETUP_negedge_posedge, `FD2TQHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `FD2TQHS_TI_CP_SETUP_posedge_posedge, `FD2TQHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `FD2TQHS_TI_CP_SETUP_negedge_posedge, `FD2TQHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `FD2TQHS_D_CP_SETUP_posedge_posedge,`FD2TQHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `FD2TQHS_D_CP_SETUP_negedge_posedge,`FD2TQHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD2TQHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2TQHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2TQHS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FD2TQHS_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `FD2TQHS_CD_CP_REM_posedge_posedge, Notifier);
`endif 
   endspecify
`endif


endmodule // FD2TQHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:52 and Version :1.1 //
 
//  START 
// CELL FD2TQHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD2TQHSP_CD_F_SO_F 0.1
`define FD2TQHSP_CP_R_SO_R 0.1
`define FD2TQHSP_CP_R_SO_F 0.1
`define FD2TQHSP_CD_F_Q_F 0.1
`define FD2TQHSP_CP_R_Q_R 0.1
`define FD2TQHSP_CP_R_Q_F 0.1
`define FD2TQHSP_CD_CP_REM_posedge_posedge 0.1
`define FD2TQHSP_CD_CP_REC_posedge_posedge 0.1
`define FD2TQHSP_CD_PWL 0.1
`define FD2TQHSP_CP_PWH 0.1
`define FD2TQHSP_CP_PWL 0.1
`define FD2TQHSP_D_CP_SETUP_posedge_posedge 0.1
`define FD2TQHSP_D_CP_SETUP_negedge_posedge 0.1
`define FD2TQHSP_D_CP_HOLD_posedge_posedge 0.1
`define FD2TQHSP_D_CP_HOLD_negedge_posedge 0.1
`define FD2TQHSP_TI_CP_SETUP_posedge_posedge 0.1
`define FD2TQHSP_TI_CP_SETUP_negedge_posedge 0.1
`define FD2TQHSP_TI_CP_HOLD_posedge_posedge 0.1
`define FD2TQHSP_TI_CP_HOLD_negedge_posedge 0.1
`define FD2TQHSP_TE_CP_SETUP_posedge_posedge 0.1
`define FD2TQHSP_TE_CP_SETUP_negedge_posedge 0.1
`define FD2TQHSP_TE_CP_HOLD_posedge_posedge 0.1
`define FD2TQHSP_TE_CP_HOLD_negedge_posedge 0.1

module FD2TQHSP (Q, SO, D, CP, CD, TI, TE);

   output Q;
   output SO;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);
   buf  u3 (SO, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   and  (AndCDTEX_, CD, TEX);
   and  (AndCDTE_, CD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && CD) (posedge CP => (Q +: D)) = (`FD2TQHSP_CP_R_Q_R, `FD2TQHSP_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`FD2TQHSP_CP_R_Q_R, `FD2TQHSP_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`FD2TQHSP_CP_R_Q_R, `FD2TQHSP_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`FD2TQHSP_CP_R_Q_R, `FD2TQHSP_CP_R_Q_F);
      if(!TE && CD) (posedge CP => (SO +: D)) = (`FD2TQHSP_CP_R_SO_R, `FD2TQHSP_CP_R_SO_F);
      if(TE && CD) (posedge CP => (SO +: TI)) = (`FD2TQHSP_CP_R_SO_R, `FD2TQHSP_CP_R_SO_F);
      if(!D && TI && CD) (posedge CP => (SO +: TE)) = (`FD2TQHSP_CP_R_SO_R, `FD2TQHSP_CP_R_SO_F);
      if(!TI && D && CD) (posedge CP => (SO -: TE)) = (`FD2TQHSP_CP_R_SO_R, `FD2TQHSP_CP_R_SO_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2TQHSP_CD_F_Q_F,`FD2TQHSP_CD_F_Q_F);
      (negedge CD => (SO +: 1'b0)) = (`FD2TQHSP_CD_F_SO_F,`FD2TQHSP_CD_F_SO_F);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FD2TQHSP_TE_CP_SETUP_posedge_posedge, `FD2TQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FD2TQHSP_TE_CP_SETUP_negedge_posedge, `FD2TQHSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `FD2TQHSP_TI_CP_SETUP_posedge_posedge, `FD2TQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `FD2TQHSP_TI_CP_SETUP_negedge_posedge, `FD2TQHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `FD2TQHSP_D_CP_SETUP_posedge_posedge, `FD2TQHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `FD2TQHSP_D_CP_SETUP_negedge_posedge, `FD2TQHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD2TQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2TQHSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2TQHSP_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FD2TQHSP_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `FD2TQHSP_CD_CP_REM_posedge_posedge, Notifier);

`else
  (posedge CP => (Q +: Mux21DTITE_)) = (`FD2TQHSP_CP_R_Q_R, `FD2TQHSP_CP_R_Q_F);
      (posedge CP => (SO +: Mux21DTITE_)) = (`FD2TQHSP_CP_R_SO_R, `FD2TQHSP_CP_R_SO_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2TQHSP_CD_F_Q_F,`FD2TQHSP_CD_F_Q_F);
      (negedge CD => (SO +: 1'b0)) = (`FD2TQHSP_CD_F_SO_F,`FD2TQHSP_CD_F_SO_F);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FD2TQHSP_TE_CP_SETUP_posedge_posedge, `FD2TQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FD2TQHSP_TE_CP_SETUP_negedge_posedge, `FD2TQHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `FD2TQHSP_TI_CP_SETUP_posedge_posedge, `FD2TQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `FD2TQHSP_TI_CP_SETUP_negedge_posedge, `FD2TQHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `FD2TQHSP_D_CP_SETUP_posedge_posedge,`FD2TQHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `FD2TQHSP_D_CP_SETUP_negedge_posedge,`FD2TQHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD2TQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2TQHSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2TQHSP_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FD2TQHSP_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `FD2TQHSP_CD_CP_REM_posedge_posedge, Notifier);
`endif 
   endspecify
`endif


endmodule // FD2TQHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:52 and Version :1.1 //
 
//  START 
// CELL FD2TQHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD2TQHSX4_CD_F_SO_F 0.1
`define FD2TQHSX4_CP_R_SO_R 0.1
`define FD2TQHSX4_CP_R_SO_F 0.1
`define FD2TQHSX4_CD_F_Q_F 0.1
`define FD2TQHSX4_CP_R_Q_R 0.1
`define FD2TQHSX4_CP_R_Q_F 0.1
`define FD2TQHSX4_CD_CP_REM_posedge_posedge 0.1
`define FD2TQHSX4_CD_CP_REC_posedge_posedge 0.1
`define FD2TQHSX4_CD_PWL 0.1
`define FD2TQHSX4_CP_PWH 0.1
`define FD2TQHSX4_CP_PWL 0.1
`define FD2TQHSX4_D_CP_SETUP_posedge_posedge 0.1
`define FD2TQHSX4_D_CP_SETUP_negedge_posedge 0.1
`define FD2TQHSX4_D_CP_HOLD_posedge_posedge 0.1
`define FD2TQHSX4_D_CP_HOLD_negedge_posedge 0.1
`define FD2TQHSX4_TI_CP_SETUP_posedge_posedge 0.1
`define FD2TQHSX4_TI_CP_SETUP_negedge_posedge 0.1
`define FD2TQHSX4_TI_CP_HOLD_posedge_posedge 0.1
`define FD2TQHSX4_TI_CP_HOLD_negedge_posedge 0.1
`define FD2TQHSX4_TE_CP_SETUP_posedge_posedge 0.1
`define FD2TQHSX4_TE_CP_SETUP_negedge_posedge 0.1
`define FD2TQHSX4_TE_CP_HOLD_posedge_posedge 0.1
`define FD2TQHSX4_TE_CP_HOLD_negedge_posedge 0.1

module FD2TQHSX4 (Q, SO, D, CP, CD, TI, TE);

   output Q;
   output SO;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);
   buf  u3 (SO, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   and  (AndCDTEX_, CD, TEX);
   and  (AndCDTE_, CD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && CD) (posedge CP => (Q +: D)) = (`FD2TQHSX4_CP_R_Q_R, `FD2TQHSX4_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`FD2TQHSX4_CP_R_Q_R, `FD2TQHSX4_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`FD2TQHSX4_CP_R_Q_R, `FD2TQHSX4_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`FD2TQHSX4_CP_R_Q_R, `FD2TQHSX4_CP_R_Q_F);
      if(!TE && CD) (posedge CP => (SO +: D)) = (`FD2TQHSX4_CP_R_SO_R, `FD2TQHSX4_CP_R_SO_F);
      if(TE && CD) (posedge CP => (SO +: TI)) = (`FD2TQHSX4_CP_R_SO_R, `FD2TQHSX4_CP_R_SO_F);
      if(!D && TI && CD) (posedge CP => (SO +: TE)) = (`FD2TQHSX4_CP_R_SO_R, `FD2TQHSX4_CP_R_SO_F);
      if(!TI && D && CD) (posedge CP => (SO -: TE)) = (`FD2TQHSX4_CP_R_SO_R, `FD2TQHSX4_CP_R_SO_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2TQHSX4_CD_F_Q_F,`FD2TQHSX4_CD_F_Q_F);
      (negedge CD => (SO +: 1'b0)) = (`FD2TQHSX4_CD_F_SO_F,`FD2TQHSX4_CD_F_SO_F);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FD2TQHSX4_TE_CP_SETUP_posedge_posedge, `FD2TQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FD2TQHSX4_TE_CP_SETUP_negedge_posedge, `FD2TQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `FD2TQHSX4_TI_CP_SETUP_posedge_posedge, `FD2TQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `FD2TQHSX4_TI_CP_SETUP_negedge_posedge, `FD2TQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `FD2TQHSX4_D_CP_SETUP_posedge_posedge, `FD2TQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `FD2TQHSX4_D_CP_SETUP_negedge_posedge, `FD2TQHSX4_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD2TQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2TQHSX4_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2TQHSX4_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FD2TQHSX4_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `FD2TQHSX4_CD_CP_REM_posedge_posedge, Notifier);

`else
  (posedge CP => (Q +: Mux21DTITE_)) = (`FD2TQHSX4_CP_R_Q_R, `FD2TQHSX4_CP_R_Q_F);
      (posedge CP => (SO +: Mux21DTITE_)) = (`FD2TQHSX4_CP_R_SO_R, `FD2TQHSX4_CP_R_SO_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2TQHSX4_CD_F_Q_F,`FD2TQHSX4_CD_F_Q_F);
      (negedge CD => (SO +: 1'b0)) = (`FD2TQHSX4_CD_F_SO_F,`FD2TQHSX4_CD_F_SO_F);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FD2TQHSX4_TE_CP_SETUP_posedge_posedge, `FD2TQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FD2TQHSX4_TE_CP_SETUP_negedge_posedge, `FD2TQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `FD2TQHSX4_TI_CP_SETUP_posedge_posedge, `FD2TQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `FD2TQHSX4_TI_CP_SETUP_negedge_posedge, `FD2TQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `FD2TQHSX4_D_CP_SETUP_posedge_posedge,`FD2TQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `FD2TQHSX4_D_CP_SETUP_negedge_posedge,`FD2TQHSX4_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD2TQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2TQHSX4_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2TQHSX4_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FD2TQHSX4_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `FD2TQHSX4_CD_CP_REM_posedge_posedge, Notifier);
`endif 
   endspecify
`endif


endmodule // FD2TQHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:52 and Version :1.1 //
 
//  START 
// CELL FDH2TQHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDH2TQHSP_CD_F_SO_F 0.1
`define FDH2TQHSP_CP_R_SO_R 0.1
`define FDH2TQHSP_CP_R_SO_F 0.1
`define FDH2TQHSP_CD_F_Q_F 0.1
`define FDH2TQHSP_CP_R_Q_R 0.1
`define FDH2TQHSP_CP_R_Q_F 0.1
`define FDH2TQHSP_CD_CP_REM_posedge_posedge 0.1
`define FDH2TQHSP_CD_CP_REC_posedge_posedge 0.1
`define FDH2TQHSP_CD_PWL 0.1
`define FDH2TQHSP_CP_PWH 0.1
`define FDH2TQHSP_CP_PWL 0.1
`define FDH2TQHSP_D_CP_SETUP_posedge_posedge 0.1
`define FDH2TQHSP_D_CP_SETUP_negedge_posedge 0.1
`define FDH2TQHSP_D_CP_HOLD_posedge_posedge 0.1
`define FDH2TQHSP_D_CP_HOLD_negedge_posedge 0.1
`define FDH2TQHSP_TI_CP_SETUP_posedge_posedge 0.1
`define FDH2TQHSP_TI_CP_SETUP_negedge_posedge 0.1
`define FDH2TQHSP_TI_CP_HOLD_posedge_posedge 0.1
`define FDH2TQHSP_TI_CP_HOLD_negedge_posedge 0.1
`define FDH2TQHSP_TE_CP_SETUP_posedge_posedge 0.1
`define FDH2TQHSP_TE_CP_SETUP_negedge_posedge 0.1
`define FDH2TQHSP_TE_CP_HOLD_posedge_posedge 0.1
`define FDH2TQHSP_TE_CP_HOLD_negedge_posedge 0.1

module FDH2TQHSP (Q, SO, D, CP, CD, TI, TE);

   output Q;
   output SO;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);
   buf  u3 (SO, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   and  (AndCDTEX_, CD, TEX);
   and  (AndCDTE_, CD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && CD) (posedge CP => (Q +: D)) = (`FDH2TQHSP_CP_R_Q_R, `FDH2TQHSP_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`FDH2TQHSP_CP_R_Q_R, `FDH2TQHSP_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`FDH2TQHSP_CP_R_Q_R, `FDH2TQHSP_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`FDH2TQHSP_CP_R_Q_R, `FDH2TQHSP_CP_R_Q_F);
      if(!TE && CD) (posedge CP => (SO +: D)) = (`FDH2TQHSP_CP_R_SO_R, `FDH2TQHSP_CP_R_SO_F);
      if(TE && CD) (posedge CP => (SO +: TI)) = (`FDH2TQHSP_CP_R_SO_R, `FDH2TQHSP_CP_R_SO_F);
      if(!D && TI && CD) (posedge CP => (SO +: TE)) = (`FDH2TQHSP_CP_R_SO_R, `FDH2TQHSP_CP_R_SO_F);
      if(!TI && D && CD) (posedge CP => (SO -: TE)) = (`FDH2TQHSP_CP_R_SO_R, `FDH2TQHSP_CP_R_SO_F);
      (negedge CD => (Q +: 1'b0)) = (`FDH2TQHSP_CD_F_Q_F,`FDH2TQHSP_CD_F_Q_F);
      (negedge CD => (SO +: 1'b0)) = (`FDH2TQHSP_CD_F_SO_F,`FDH2TQHSP_CD_F_SO_F);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FDH2TQHSP_TE_CP_SETUP_posedge_posedge, `FDH2TQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FDH2TQHSP_TE_CP_SETUP_negedge_posedge, `FDH2TQHSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `FDH2TQHSP_TI_CP_SETUP_posedge_posedge, `FDH2TQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `FDH2TQHSP_TI_CP_SETUP_negedge_posedge, `FDH2TQHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `FDH2TQHSP_D_CP_SETUP_posedge_posedge, `FDH2TQHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `FDH2TQHSP_D_CP_SETUP_negedge_posedge, `FDH2TQHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDH2TQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDH2TQHSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDH2TQHSP_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FDH2TQHSP_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `FDH2TQHSP_CD_CP_REM_posedge_posedge, Notifier);

`else
  (posedge CP => (Q +: Mux21DTITE_)) = (`FDH2TQHSP_CP_R_Q_R, `FDH2TQHSP_CP_R_Q_F);
      (posedge CP => (SO +: Mux21DTITE_)) = (`FDH2TQHSP_CP_R_SO_R, `FDH2TQHSP_CP_R_SO_F);
      (negedge CD => (Q +: 1'b0)) = (`FDH2TQHSP_CD_F_Q_F,`FDH2TQHSP_CD_F_Q_F);
      (negedge CD => (SO +: 1'b0)) = (`FDH2TQHSP_CD_F_SO_F,`FDH2TQHSP_CD_F_SO_F);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FDH2TQHSP_TE_CP_SETUP_posedge_posedge, `FDH2TQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FDH2TQHSP_TE_CP_SETUP_negedge_posedge, `FDH2TQHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `FDH2TQHSP_TI_CP_SETUP_posedge_posedge, `FDH2TQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `FDH2TQHSP_TI_CP_SETUP_negedge_posedge, `FDH2TQHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `FDH2TQHSP_D_CP_SETUP_posedge_posedge,`FDH2TQHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `FDH2TQHSP_D_CP_SETUP_negedge_posedge,`FDH2TQHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDH2TQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDH2TQHSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDH2TQHSP_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FDH2TQHSP_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `FDH2TQHSP_CD_CP_REM_posedge_posedge, Notifier);
`endif 
   endspecify
`endif


endmodule // FDH2TQHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:52 and Version :1.1 //
 
//  START 
// CELL FDH2TQHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDH2TQHSX4_CD_F_SO_F 0.1
`define FDH2TQHSX4_CP_R_SO_R 0.1
`define FDH2TQHSX4_CP_R_SO_F 0.1
`define FDH2TQHSX4_CD_F_Q_F 0.1
`define FDH2TQHSX4_CP_R_Q_R 0.1
`define FDH2TQHSX4_CP_R_Q_F 0.1
`define FDH2TQHSX4_CD_CP_REM_posedge_posedge 0.1
`define FDH2TQHSX4_CD_CP_REC_posedge_posedge 0.1
`define FDH2TQHSX4_CD_PWL 0.1
`define FDH2TQHSX4_CP_PWH 0.1
`define FDH2TQHSX4_CP_PWL 0.1
`define FDH2TQHSX4_D_CP_SETUP_posedge_posedge 0.1
`define FDH2TQHSX4_D_CP_SETUP_negedge_posedge 0.1
`define FDH2TQHSX4_D_CP_HOLD_posedge_posedge 0.1
`define FDH2TQHSX4_D_CP_HOLD_negedge_posedge 0.1
`define FDH2TQHSX4_TI_CP_SETUP_posedge_posedge 0.1
`define FDH2TQHSX4_TI_CP_SETUP_negedge_posedge 0.1
`define FDH2TQHSX4_TI_CP_HOLD_posedge_posedge 0.1
`define FDH2TQHSX4_TI_CP_HOLD_negedge_posedge 0.1
`define FDH2TQHSX4_TE_CP_SETUP_posedge_posedge 0.1
`define FDH2TQHSX4_TE_CP_SETUP_negedge_posedge 0.1
`define FDH2TQHSX4_TE_CP_HOLD_posedge_posedge 0.1
`define FDH2TQHSX4_TE_CP_HOLD_negedge_posedge 0.1

module FDH2TQHSX4 (Q, SO, D, CP, CD, TI, TE);

   output Q;
   output SO;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);
   buf  u3 (SO, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   and  (AndCDTEX_, CD, TEX);
   and  (AndCDTE_, CD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && CD) (posedge CP => (Q +: D)) = (`FDH2TQHSX4_CP_R_Q_R, `FDH2TQHSX4_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`FDH2TQHSX4_CP_R_Q_R, `FDH2TQHSX4_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`FDH2TQHSX4_CP_R_Q_R, `FDH2TQHSX4_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`FDH2TQHSX4_CP_R_Q_R, `FDH2TQHSX4_CP_R_Q_F);
      if(!TE && CD) (posedge CP => (SO +: D)) = (`FDH2TQHSX4_CP_R_SO_R, `FDH2TQHSX4_CP_R_SO_F);
      if(TE && CD) (posedge CP => (SO +: TI)) = (`FDH2TQHSX4_CP_R_SO_R, `FDH2TQHSX4_CP_R_SO_F);
      if(!D && TI && CD) (posedge CP => (SO +: TE)) = (`FDH2TQHSX4_CP_R_SO_R, `FDH2TQHSX4_CP_R_SO_F);
      if(!TI && D && CD) (posedge CP => (SO -: TE)) = (`FDH2TQHSX4_CP_R_SO_R, `FDH2TQHSX4_CP_R_SO_F);
      (negedge CD => (Q +: 1'b0)) = (`FDH2TQHSX4_CD_F_Q_F,`FDH2TQHSX4_CD_F_Q_F);
      (negedge CD => (SO +: 1'b0)) = (`FDH2TQHSX4_CD_F_SO_F,`FDH2TQHSX4_CD_F_SO_F);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FDH2TQHSX4_TE_CP_SETUP_posedge_posedge, `FDH2TQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FDH2TQHSX4_TE_CP_SETUP_negedge_posedge, `FDH2TQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `FDH2TQHSX4_TI_CP_SETUP_posedge_posedge, `FDH2TQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `FDH2TQHSX4_TI_CP_SETUP_negedge_posedge, `FDH2TQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `FDH2TQHSX4_D_CP_SETUP_posedge_posedge, `FDH2TQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `FDH2TQHSX4_D_CP_SETUP_negedge_posedge, `FDH2TQHSX4_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDH2TQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDH2TQHSX4_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDH2TQHSX4_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FDH2TQHSX4_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `FDH2TQHSX4_CD_CP_REM_posedge_posedge, Notifier);

`else
  (posedge CP => (Q +: Mux21DTITE_)) = (`FDH2TQHSX4_CP_R_Q_R, `FDH2TQHSX4_CP_R_Q_F);
      (posedge CP => (SO +: Mux21DTITE_)) = (`FDH2TQHSX4_CP_R_SO_R, `FDH2TQHSX4_CP_R_SO_F);
      (negedge CD => (Q +: 1'b0)) = (`FDH2TQHSX4_CD_F_Q_F,`FDH2TQHSX4_CD_F_Q_F);
      (negedge CD => (SO +: 1'b0)) = (`FDH2TQHSX4_CD_F_SO_F,`FDH2TQHSX4_CD_F_SO_F);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FDH2TQHSX4_TE_CP_SETUP_posedge_posedge, `FDH2TQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FDH2TQHSX4_TE_CP_SETUP_negedge_posedge, `FDH2TQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `FDH2TQHSX4_TI_CP_SETUP_posedge_posedge, `FDH2TQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `FDH2TQHSX4_TI_CP_SETUP_negedge_posedge, `FDH2TQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `FDH2TQHSX4_D_CP_SETUP_posedge_posedge,`FDH2TQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `FDH2TQHSX4_D_CP_SETUP_negedge_posedge,`FDH2TQHSX4_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDH2TQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDH2TQHSX4_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDH2TQHSX4_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FDH2TQHSX4_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `FDH2TQHSX4_CD_CP_REM_posedge_posedge, Notifier);
`endif 
   endspecify
`endif


endmodule // FDH2TQHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:52 and Version :1.1 //
 
//  START 
// CELL FDH2TQHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDH2TQHSX8_CD_F_SO_F 0.1
`define FDH2TQHSX8_CP_R_SO_R 0.1
`define FDH2TQHSX8_CP_R_SO_F 0.1
`define FDH2TQHSX8_CD_F_Q_F 0.1
`define FDH2TQHSX8_CP_R_Q_R 0.1
`define FDH2TQHSX8_CP_R_Q_F 0.1
`define FDH2TQHSX8_CD_CP_REM_posedge_posedge 0.1
`define FDH2TQHSX8_CD_CP_REC_posedge_posedge 0.1
`define FDH2TQHSX8_CD_PWL 0.1
`define FDH2TQHSX8_CP_PWH 0.1
`define FDH2TQHSX8_CP_PWL 0.1
`define FDH2TQHSX8_D_CP_SETUP_posedge_posedge 0.1
`define FDH2TQHSX8_D_CP_SETUP_negedge_posedge 0.1
`define FDH2TQHSX8_D_CP_HOLD_posedge_posedge 0.1
`define FDH2TQHSX8_D_CP_HOLD_negedge_posedge 0.1
`define FDH2TQHSX8_TI_CP_SETUP_posedge_posedge 0.1
`define FDH2TQHSX8_TI_CP_SETUP_negedge_posedge 0.1
`define FDH2TQHSX8_TI_CP_HOLD_posedge_posedge 0.1
`define FDH2TQHSX8_TI_CP_HOLD_negedge_posedge 0.1
`define FDH2TQHSX8_TE_CP_SETUP_posedge_posedge 0.1
`define FDH2TQHSX8_TE_CP_SETUP_negedge_posedge 0.1
`define FDH2TQHSX8_TE_CP_HOLD_posedge_posedge 0.1
`define FDH2TQHSX8_TE_CP_HOLD_negedge_posedge 0.1

module FDH2TQHSX8 (Q, SO, D, CP, CD, TI, TE);

   output Q;
   output SO;
   input D;
   input CP;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2 u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, Notifier);

   buf  u2 (Q, IQ);
   buf  u3 (SO, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   and  (AndCDTEX_, CD, TEX);
   and  (AndCDTE_, CD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && CD) (posedge CP => (Q +: D)) = (`FDH2TQHSX8_CP_R_Q_R, `FDH2TQHSX8_CP_R_Q_F);
      if(TE && CD) (posedge CP => (Q +: TI)) = (`FDH2TQHSX8_CP_R_Q_R, `FDH2TQHSX8_CP_R_Q_F);
      if(!D && TI && CD) (posedge CP => (Q +: TE)) = (`FDH2TQHSX8_CP_R_Q_R, `FDH2TQHSX8_CP_R_Q_F);
      if(!TI && D && CD) (posedge CP => (Q -: TE)) = (`FDH2TQHSX8_CP_R_Q_R, `FDH2TQHSX8_CP_R_Q_F);
      if(!TE && CD) (posedge CP => (SO +: D)) = (`FDH2TQHSX8_CP_R_SO_R, `FDH2TQHSX8_CP_R_SO_F);
      if(TE && CD) (posedge CP => (SO +: TI)) = (`FDH2TQHSX8_CP_R_SO_R, `FDH2TQHSX8_CP_R_SO_F);
      if(!D && TI && CD) (posedge CP => (SO +: TE)) = (`FDH2TQHSX8_CP_R_SO_R, `FDH2TQHSX8_CP_R_SO_F);
      if(!TI && D && CD) (posedge CP => (SO -: TE)) = (`FDH2TQHSX8_CP_R_SO_R, `FDH2TQHSX8_CP_R_SO_F);
      (negedge CD => (Q +: 1'b0)) = (`FDH2TQHSX8_CD_F_Q_F,`FDH2TQHSX8_CD_F_Q_F);
      (negedge CD => (SO +: 1'b0)) = (`FDH2TQHSX8_CD_F_SO_F,`FDH2TQHSX8_CD_F_SO_F);

	$setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FDH2TQHSX8_TE_CP_SETUP_posedge_posedge, `FDH2TQHSX8_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FDH2TQHSX8_TE_CP_SETUP_negedge_posedge, `FDH2TQHSX8_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTE_, posedge TI, `FDH2TQHSX8_TI_CP_SETUP_posedge_posedge, `FDH2TQHSX8_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTE_, negedge TI, `FDH2TQHSX8_TI_CP_SETUP_negedge_posedge, `FDH2TQHSX8_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDTEX_, posedge D, `FDH2TQHSX8_D_CP_SETUP_posedge_posedge, `FDH2TQHSX8_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDTEX_, negedge D, `FDH2TQHSX8_D_CP_SETUP_negedge_posedge, `FDH2TQHSX8_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDH2TQHSX8_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDH2TQHSX8_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDH2TQHSX8_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FDH2TQHSX8_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& Mux21DTITE_, posedge CD, `FDH2TQHSX8_CD_CP_REM_posedge_posedge, Notifier);

`else
  (posedge CP => (Q +: Mux21DTITE_)) = (`FDH2TQHSX8_CP_R_Q_R, `FDH2TQHSX8_CP_R_Q_F);
      (posedge CP => (SO +: Mux21DTITE_)) = (`FDH2TQHSX8_CP_R_SO_R, `FDH2TQHSX8_CP_R_SO_F);
      (negedge CD => (Q +: 1'b0)) = (`FDH2TQHSX8_CD_F_Q_F,`FDH2TQHSX8_CD_F_Q_F);
      (negedge CD => (SO +: 1'b0)) = (`FDH2TQHSX8_CD_F_SO_F,`FDH2TQHSX8_CD_F_SO_F);
 
        $setuphold(posedge CP &&& AndXorDTI_CD_, posedge TE, `FDH2TQHSX8_TE_CP_SETUP_posedge_posedge, `FDH2TQHSX8_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CD_, negedge TE, `FDH2TQHSX8_TE_CP_SETUP_negedge_posedge, `FDH2TQHSX8_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTE_, posedge TI, `FDH2TQHSX8_TI_CP_SETUP_posedge_posedge, `FDH2TQHSX8_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTE_, negedge TI, `FDH2TQHSX8_TI_CP_SETUP_negedge_posedge, `FDH2TQHSX8_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDTEX_, posedge D, `FDH2TQHSX8_D_CP_SETUP_posedge_posedge,`FDH2TQHSX8_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDTEX_, negedge D, `FDH2TQHSX8_D_CP_SETUP_negedge_posedge,`FDH2TQHSX8_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDH2TQHSX8_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FDH2TQHSX8_CP_PWH, 0, Notifier);
      $width(negedge CD, `FDH2TQHSX8_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& Mux21DTITE_, `FDH2TQHSX8_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& Mux21DTITE_, posedge CD, `FDH2TQHSX8_CD_CP_REM_posedge_posedge, Notifier);
`endif 
   endspecify
`endif


endmodule // FDH2TQHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:52 and Version :1.1 //
 
//  START 
// CELL FD2_SYNCHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD2_SYNCHS_CD_F_QN_R 0.1
`define FD2_SYNCHS_CP_R_QN_F 0.1
`define FD2_SYNCHS_CP_R_QN_R 0.1
`define FD2_SYNCHS_CD_F_Q_F 0.1
`define FD2_SYNCHS_CP_R_Q_R 0.1
`define FD2_SYNCHS_CP_R_Q_F 0.1
`define FD2_SYNCHS_CD_CP_REM_posedge_posedge 0.1
`define FD2_SYNCHS_CD_CP_REC_posedge_posedge 0.1
`define FD2_SYNCHS_CD_PWL 0.1
`define FD2_SYNCHS_CP_PWH 0.1
`define FD2_SYNCHS_CP_PWL 0.1
`define FD2_SYNCHS_D_CP_SETUP_posedge_posedge 0.1
`define FD2_SYNCHS_D_CP_SETUP_negedge_posedge 0.1
`define FD2_SYNCHS_D_CP_HOLD_posedge_posedge 0.1
`define FD2_SYNCHS_D_CP_HOLD_negedge_posedge 0.1

module FD2_SYNCHS (Q, QN, D, CP, CD);

   output Q;
   output QN;
   input D;
   input CP;
   input CD;


   reg Notifier;


   U_FD_P_RN_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, CD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   specify
`ifdef verifault
      if(CD) (posedge CP => (Q +: D)) = (`FD2_SYNCHS_CP_R_Q_R, `FD2_SYNCHS_CP_R_Q_F);
      if(CD) (posedge CP => (QN -: D)) = (`FD2_SYNCHS_CP_R_QN_R, `FD2_SYNCHS_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2_SYNCHS_CD_F_Q_F,`FD2_SYNCHS_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FD2_SYNCHS_CD_F_QN_R,`FD2_SYNCHS_CD_F_QN_R);

	$setuphold(posedge CP &&& CD, posedge D, `FD2_SYNCHS_D_CP_SETUP_posedge_posedge, `FD2_SYNCHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge D, `FD2_SYNCHS_D_CP_SETUP_negedge_posedge, `FD2_SYNCHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD2_SYNCHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2_SYNCHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2_SYNCHS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& D, `FD2_SYNCHS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D, posedge CD, `FD2_SYNCHS_CD_CP_REM_posedge_posedge, Notifier);
`else

      (posedge CP => (Q +: D)) = (`FD2_SYNCHS_CP_R_Q_R, `FD2_SYNCHS_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`FD2_SYNCHS_CP_R_QN_R, `FD2_SYNCHS_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FD2_SYNCHS_CD_F_Q_F,`FD2_SYNCHS_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FD2_SYNCHS_CD_F_QN_R,`FD2_SYNCHS_CD_F_QN_R);
 
        $setuphold(posedge CP &&& CD, posedge D, `FD2_SYNCHS_D_CP_SETUP_posedge_posedge, `FD2_SYNCHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge D, `FD2_SYNCHS_D_CP_SETUP_negedge_posedge, `FD2_SYNCHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD2_SYNCHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FD2_SYNCHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FD2_SYNCHS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& D, `FD2_SYNCHS_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D, posedge CD, `FD2_SYNCHS_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FD2_SYNCHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:20 and Version :1.1 //
 
//  START 
// CELL FD3HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD3HS_SD_F_QN_F 0.1
`define FD3HS_CD_F_QN_R 0.1
`define FD3HS_CD_R_QN_F 0.1
`define FD3HS_CP_R_QN_F 0.1
`define FD3HS_CP_R_QN_R 0.1
`define FD3HS_SD_F_Q_R 0.1
`define FD3HS_CD_F_Q_F 0.1
`define FD3HS_CD_R_Q_R 0.1
`define FD3HS_CP_R_Q_R 0.1
`define FD3HS_CP_R_Q_F 0.1
`define FD3HS_CD_SD_REM_posedge_posedge 0.1
`define FD3HS_CD_SD_REC_posedge_posedge 0.1
`define FD3HS_CD_CP_REM_posedge_posedge 0.1
`define FD3HS_SD_CP_REM_posedge_posedge 0.1
`define FD3HS_CD_CP_REC_posedge_posedge 0.1
`define FD3HS_SD_CP_REC_posedge_posedge 0.1
`define FD3HS_CD_PWL 0.1
`define FD3HS_SD_PWL 0.1
`define FD3HS_CP_PWH 0.1
`define FD3HS_CP_PWL 0.1
`define FD3HS_D_CP_SETUP_posedge_posedge 0.1
`define FD3HS_D_CP_SETUP_negedge_posedge 0.1
`define FD3HS_D_CP_HOLD_posedge_posedge 0.1
`define FD3HS_D_CP_HOLD_negedge_posedge 0.1

module FD3HS (Q, QN, D, CP, CD, SD);

   output Q;
   output QN;
   input D;
   input CP;
   input CD;
   input SD;


   reg Notifier;


   U_FD_P_RN_SN_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, CD, SD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);




`ifdef functional
`else
   and  (AndCDSD_, CD, SD);
 
   and  (AndSDD, SD, D);
   not  (D_, D);
   and  (AndCDD_, CD, D_);

   specify
`ifdef verifault

      if(CD && SD) (posedge CP => (Q +: D)) = (`FD3HS_CP_R_Q_R, `FD3HS_CP_R_Q_F);
      if(CD && SD) (posedge CP => (QN -: D)) = (`FD3HS_CP_R_QN_R, `FD3HS_CP_R_QN_F);
      if(!SD) (posedge CD => (Q +: 1'b1)) = (`FD3HS_CD_R_Q_R,`FD3HS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3HS_CD_R_Q_R,`FD3HS_CD_F_Q_F);
      if(CD) (negedge SD => (Q +: 1'b1)) = (`FD3HS_SD_F_Q_R,`FD3HS_SD_F_Q_R);
      if(!SD) (posedge CD => (QN +: 1'b0)) = (`FD3HS_CD_F_QN_R,`FD3HS_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`FD3HS_CD_F_QN_R,`FD3HS_CD_R_QN_F);
      if(CD) (negedge SD => (QN +: 1'b0)) = (`FD3HS_SD_F_QN_F,`FD3HS_SD_F_QN_F);

	$setuphold(posedge CP &&& AndCDSD_, posedge D, `FD3HS_D_CP_SETUP_posedge_posedge, `FD3HS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSD_, negedge D, `FD3HS_D_CP_SETUP_negedge_posedge, `FD3HS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD3HS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3HS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3HS_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3HS_CD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& AndCDD_, `FD3HS_SD_CP_REC_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge CP &&& AndSDD, `FD3HS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndCDD_, posedge SD, `FD3HS_SD_CP_REM_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndSDD, posedge CD, `FD3HS_CD_CP_REM_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge SD, `FD3HS_CD_SD_REC_posedge_posedge, Notifier);

	$hold(posedge SD, posedge CD, `FD3HS_CD_SD_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: D)) = (`FD3HS_CP_R_Q_R, `FD3HS_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`FD3HS_CP_R_QN_R, `FD3HS_CP_R_QN_F);
      (posedge CD => (Q +: 1'b1)) = (`FD3HS_CD_R_Q_R,`FD3HS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3HS_CD_R_Q_R,`FD3HS_CD_F_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD3HS_SD_F_Q_R,`FD3HS_SD_F_Q_R);
      (posedge CD => (QN +: 1'b0)) = (`FD3HS_CD_F_QN_R,`FD3HS_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`FD3HS_CD_F_QN_R,`FD3HS_CD_R_QN_F);
      (negedge SD => (QN +: 1'b0)) = (`FD3HS_SD_F_QN_F,`FD3HS_SD_F_QN_F);
 
        $setuphold(posedge CP &&& AndCDSD_, posedge D, `FD3HS_D_CP_SETUP_posedge_posedge, `FD3HS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSD_, negedge D, `FD3HS_D_CP_SETUP_negedge_posedge, `FD3HS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD3HS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3HS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3HS_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3HS_CD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& AndCDD_, `FD3HS_SD_CP_REC_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge CP &&& AndSDD, `FD3HS_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndCDD_, posedge SD, `FD3HS_SD_CP_REM_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndSDD, posedge CD, `FD3HS_CD_CP_REM_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge SD, `FD3HS_CD_SD_REC_posedge_posedge, Notifier);
        $hold(posedge SD, posedge CD, `FD3HS_CD_SD_REM_posedge_posedge, Notifier);

`endif
   endspecify
`endif

endmodule // FD3HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:58 and Version :1.1 //
 
//  START 
// CELL FD3HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD3HSP_SD_F_QN_F 0.1
`define FD3HSP_CD_F_QN_R 0.1
`define FD3HSP_CD_R_QN_F 0.1
`define FD3HSP_CP_R_QN_F 0.1
`define FD3HSP_CP_R_QN_R 0.1
`define FD3HSP_SD_F_Q_R 0.1
`define FD3HSP_CD_F_Q_F 0.1
`define FD3HSP_CD_R_Q_R 0.1
`define FD3HSP_CP_R_Q_R 0.1
`define FD3HSP_CP_R_Q_F 0.1
`define FD3HSP_CD_SD_REM_posedge_posedge 0.1
`define FD3HSP_CD_SD_REC_posedge_posedge 0.1
`define FD3HSP_CD_CP_REM_posedge_posedge 0.1
`define FD3HSP_SD_CP_REM_posedge_posedge 0.1
`define FD3HSP_CD_CP_REC_posedge_posedge 0.1
`define FD3HSP_SD_CP_REC_posedge_posedge 0.1
`define FD3HSP_CD_PWL 0.1
`define FD3HSP_SD_PWL 0.1
`define FD3HSP_CP_PWH 0.1
`define FD3HSP_CP_PWL 0.1
`define FD3HSP_D_CP_SETUP_posedge_posedge 0.1
`define FD3HSP_D_CP_SETUP_negedge_posedge 0.1
`define FD3HSP_D_CP_HOLD_posedge_posedge 0.1
`define FD3HSP_D_CP_HOLD_negedge_posedge 0.1

module FD3HSP (Q, QN, D, CP, CD, SD);

   output Q;
   output QN;
   input D;
   input CP;
   input CD;
   input SD;


   reg Notifier;


   U_FD_P_RN_SN_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, CD, SD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);




`ifdef functional
`else
   and  (AndCDSD_, CD, SD);
 
   and  (AndSDD, SD, D);
   not  (D_, D);
   and  (AndCDD_, CD, D_);

   specify
`ifdef verifault

      if(CD && SD) (posedge CP => (Q +: D)) = (`FD3HSP_CP_R_Q_R, `FD3HSP_CP_R_Q_F);
      if(CD && SD) (posedge CP => (QN -: D)) = (`FD3HSP_CP_R_QN_R, `FD3HSP_CP_R_QN_F);
      if(!SD) (posedge CD => (Q +: 1'b1)) = (`FD3HSP_CD_R_Q_R,`FD3HSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3HSP_CD_R_Q_R,`FD3HSP_CD_F_Q_F);
      if(CD) (negedge SD => (Q +: 1'b1)) = (`FD3HSP_SD_F_Q_R,`FD3HSP_SD_F_Q_R);
      if(!SD) (posedge CD => (QN +: 1'b0)) = (`FD3HSP_CD_F_QN_R,`FD3HSP_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`FD3HSP_CD_F_QN_R,`FD3HSP_CD_R_QN_F);
      if(CD) (negedge SD => (QN +: 1'b0)) = (`FD3HSP_SD_F_QN_F,`FD3HSP_SD_F_QN_F);

	$setuphold(posedge CP &&& AndCDSD_, posedge D, `FD3HSP_D_CP_SETUP_posedge_posedge, `FD3HSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSD_, negedge D, `FD3HSP_D_CP_SETUP_negedge_posedge, `FD3HSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD3HSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3HSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3HSP_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3HSP_CD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& AndCDD_, `FD3HSP_SD_CP_REC_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge CP &&& AndSDD, `FD3HSP_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndCDD_, posedge SD, `FD3HSP_SD_CP_REM_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndSDD, posedge CD, `FD3HSP_CD_CP_REM_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge SD, `FD3HSP_CD_SD_REC_posedge_posedge, Notifier);

	$hold(posedge SD, posedge CD, `FD3HSP_CD_SD_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: D)) = (`FD3HSP_CP_R_Q_R, `FD3HSP_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`FD3HSP_CP_R_QN_R, `FD3HSP_CP_R_QN_F);
      (posedge CD => (Q +: 1'b1)) = (`FD3HSP_CD_R_Q_R,`FD3HSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3HSP_CD_R_Q_R,`FD3HSP_CD_F_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD3HSP_SD_F_Q_R,`FD3HSP_SD_F_Q_R);
      (posedge CD => (QN +: 1'b0)) = (`FD3HSP_CD_F_QN_R,`FD3HSP_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`FD3HSP_CD_F_QN_R,`FD3HSP_CD_R_QN_F);
      (negedge SD => (QN +: 1'b0)) = (`FD3HSP_SD_F_QN_F,`FD3HSP_SD_F_QN_F);
 
        $setuphold(posedge CP &&& AndCDSD_, posedge D, `FD3HSP_D_CP_SETUP_posedge_posedge, `FD3HSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSD_, negedge D, `FD3HSP_D_CP_SETUP_negedge_posedge, `FD3HSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD3HSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3HSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3HSP_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3HSP_CD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& AndCDD_, `FD3HSP_SD_CP_REC_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge CP &&& AndSDD, `FD3HSP_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndCDD_, posedge SD, `FD3HSP_SD_CP_REM_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndSDD, posedge CD, `FD3HSP_CD_CP_REM_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge SD, `FD3HSP_CD_SD_REC_posedge_posedge, Notifier);
        $hold(posedge SD, posedge CD, `FD3HSP_CD_SD_REM_posedge_posedge, Notifier);

`endif
   endspecify
`endif

endmodule // FD3HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:15:58 and Version :1.1 //
 
//  START 
// CELL FD3QHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD3QHS_SD_F_Q_R 0.1
`define FD3QHS_CD_F_Q_F 0.1
`define FD3QHS_CD_R_Q_R 0.1
`define FD3QHS_CP_R_Q_R 0.1
`define FD3QHS_CP_R_Q_F 0.1
`define FD3QHS_D_CP_HOLD_posedge_posedge 0.1
`define FD3QHS_D_CP_HOLD_negedge_posedge 0.1
`define FD3QHS_D_CP_SETUP_posedge_posedge 0.1
`define FD3QHS_D_CP_SETUP_negedge_posedge 0.1
`define FD3QHS_CP_PWL 0.1
`define FD3QHS_CP_PWH 0.1
`define FD3QHS_SD_PWL 0.1
`define FD3QHS_CD_PWL 0.1
`define FD3QHS_SD_CP_REC_posedge_posedge 0.1
`define FD3QHS_CD_CP_REC_posedge_posedge 0.1
`define FD3QHS_SD_CP_REM_posedge_posedge 0.1
`define FD3QHS_CD_CP_REM_posedge_posedge 0.1
`define FD3QHS_CD_SD_REC_posedge_posedge 0.1
`define FD3QHS_CD_SD_REM_posedge_posedge 0.1

module FD3QHS (Q, D, CP, CD, SD);

   output Q;
   input D;
   input CP;
   input CD;
   input SD;


   reg Notifier;


   U_FD_P_RN_SN_NOTI u0 (IQ, D, CP, CD, SD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   and  (AndCDSD_, CD, SD);
 
   and  (AndSDD, SD, D);
   not  (D_, D);
   and  (AndCDD_, CD, D_);

   specify
`ifdef verifault

      if(CD && SD) (posedge CP => (Q +: D)) = (`FD3QHS_CP_R_Q_R, `FD3QHS_CP_R_Q_F);
      if(!SD) (posedge CD => (Q +: 1'b1)) = (`FD3QHS_CD_R_Q_R,`FD3QHS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3QHS_CD_R_Q_R,`FD3QHS_CD_F_Q_F);
      if(CD) (negedge SD => (Q +: 1'b1)) = (`FD3QHS_SD_F_Q_R,`FD3QHS_SD_F_Q_R);

	$setuphold(posedge CP &&& AndCDSD_, posedge D, `FD3QHS_D_CP_SETUP_posedge_posedge, `FD3QHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSD_, negedge D, `FD3QHS_D_CP_SETUP_negedge_posedge, `FD3QHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD3QHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3QHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3QHS_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3QHS_CD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& AndCDD_, `FD3QHS_SD_CP_REC_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge CP &&& AndSDD, `FD3QHS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndCDD_, posedge SD, `FD3QHS_SD_CP_REM_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndSDD, posedge CD, `FD3QHS_CD_CP_REM_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge SD, `FD3QHS_CD_SD_REC_posedge_posedge, Notifier);

	$hold(posedge SD, posedge CD, `FD3QHS_CD_SD_REM_posedge_posedge, Notifier);
`else
      (posedge CP => (Q +: D)) = (`FD3QHS_CP_R_Q_R, `FD3QHS_CP_R_Q_F);
      (posedge CD => (Q +: 1'b1)) = (`FD3QHS_CD_R_Q_R,`FD3QHS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3QHS_CD_R_Q_R,`FD3QHS_CD_F_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD3QHS_SD_F_Q_R,`FD3QHS_SD_F_Q_R);
 
        $setuphold(posedge CP &&& AndCDSD_, posedge D, `FD3QHS_D_CP_SETUP_posedge_posedge, `FD3QHS_D_CP_HOLD_posedge_posedge, Notifier);
 $setuphold(posedge CP &&& AndCDSD_, negedge D, `FD3QHS_D_CP_SETUP_negedge_posedge, `FD3QHS_D_CP_HOLD_negedge_posedge, Notifier);
      $width(negedge CP, `FD3QHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3QHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3QHS_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3QHS_CD_PWL, 0, Notifier);
      $recovery(posedge SD, posedge CP &&& AndCDD_, `FD3QHS_SD_CP_REC_posedge_posedge, Notifier);
 
   $recovery(posedge CD, posedge CP &&& AndSDD, `FD3QHS_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndCDD_, posedge SD, `FD3QHS_SD_CP_REM_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndSDD, posedge CD, `FD3QHS_CD_CP_REM_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge SD, `FD3QHS_CD_SD_REC_posedge_posedge, Notifier);
 
        $hold(posedge SD, posedge CD, `FD3QHS_CD_SD_REM_posedge_posedge, Notifier);
 
 
`endif

   endspecify
`endif


endmodule // FD3QHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:02 and Version :1.1 //
 
//  START 
// CELL FD3QHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD3QHSP_SD_F_Q_R 0.1
`define FD3QHSP_CD_F_Q_F 0.1
`define FD3QHSP_CD_R_Q_R 0.1
`define FD3QHSP_CP_R_Q_R 0.1
`define FD3QHSP_CP_R_Q_F 0.1
`define FD3QHSP_D_CP_HOLD_posedge_posedge 0.1
`define FD3QHSP_D_CP_HOLD_negedge_posedge 0.1
`define FD3QHSP_D_CP_SETUP_posedge_posedge 0.1
`define FD3QHSP_D_CP_SETUP_negedge_posedge 0.1
`define FD3QHSP_CP_PWL 0.1
`define FD3QHSP_CP_PWH 0.1
`define FD3QHSP_SD_PWL 0.1
`define FD3QHSP_CD_PWL 0.1
`define FD3QHSP_SD_CP_REC_posedge_posedge 0.1
`define FD3QHSP_CD_CP_REC_posedge_posedge 0.1
`define FD3QHSP_SD_CP_REM_posedge_posedge 0.1
`define FD3QHSP_CD_CP_REM_posedge_posedge 0.1
`define FD3QHSP_CD_SD_REC_posedge_posedge 0.1
`define FD3QHSP_CD_SD_REM_posedge_posedge 0.1

module FD3QHSP (Q, D, CP, CD, SD);

   output Q;
   input D;
   input CP;
   input CD;
   input SD;


   reg Notifier;


   U_FD_P_RN_SN_NOTI u0 (IQ, D, CP, CD, SD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   and  (AndCDSD_, CD, SD);
 
   and  (AndSDD, SD, D);
   not  (D_, D);
   and  (AndCDD_, CD, D_);

   specify
`ifdef verifault

      if(CD && SD) (posedge CP => (Q +: D)) = (`FD3QHSP_CP_R_Q_R, `FD3QHSP_CP_R_Q_F);
      if(!SD) (posedge CD => (Q +: 1'b1)) = (`FD3QHSP_CD_R_Q_R,`FD3QHSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3QHSP_CD_R_Q_R,`FD3QHSP_CD_F_Q_F);
      if(CD) (negedge SD => (Q +: 1'b1)) = (`FD3QHSP_SD_F_Q_R,`FD3QHSP_SD_F_Q_R);

	$setuphold(posedge CP &&& AndCDSD_, posedge D, `FD3QHSP_D_CP_SETUP_posedge_posedge, `FD3QHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSD_, negedge D, `FD3QHSP_D_CP_SETUP_negedge_posedge, `FD3QHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD3QHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3QHSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3QHSP_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3QHSP_CD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& AndCDD_, `FD3QHSP_SD_CP_REC_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge CP &&& AndSDD, `FD3QHSP_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndCDD_, posedge SD, `FD3QHSP_SD_CP_REM_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndSDD, posedge CD, `FD3QHSP_CD_CP_REM_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge SD, `FD3QHSP_CD_SD_REC_posedge_posedge, Notifier);

	$hold(posedge SD, posedge CD, `FD3QHSP_CD_SD_REM_posedge_posedge, Notifier);
`else
      (posedge CP => (Q +: D)) = (`FD3QHSP_CP_R_Q_R, `FD3QHSP_CP_R_Q_F);
      (posedge CD => (Q +: 1'b1)) = (`FD3QHSP_CD_R_Q_R,`FD3QHSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3QHSP_CD_R_Q_R,`FD3QHSP_CD_F_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD3QHSP_SD_F_Q_R,`FD3QHSP_SD_F_Q_R);
 
        $setuphold(posedge CP &&& AndCDSD_, posedge D, `FD3QHSP_D_CP_SETUP_posedge_posedge, `FD3QHSP_D_CP_HOLD_posedge_posedge, Notifier);
 $setuphold(posedge CP &&& AndCDSD_, negedge D, `FD3QHSP_D_CP_SETUP_negedge_posedge, `FD3QHSP_D_CP_HOLD_negedge_posedge, Notifier);
      $width(negedge CP, `FD3QHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3QHSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3QHSP_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3QHSP_CD_PWL, 0, Notifier);
      $recovery(posedge SD, posedge CP &&& AndCDD_, `FD3QHSP_SD_CP_REC_posedge_posedge, Notifier);
 
   $recovery(posedge CD, posedge CP &&& AndSDD, `FD3QHSP_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndCDD_, posedge SD, `FD3QHSP_SD_CP_REM_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndSDD, posedge CD, `FD3QHSP_CD_CP_REM_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge SD, `FD3QHSP_CD_SD_REC_posedge_posedge, Notifier);
 
        $hold(posedge SD, posedge CD, `FD3QHSP_CD_SD_REM_posedge_posedge, Notifier);
 
 
`endif

   endspecify
`endif


endmodule // FD3QHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:02 and Version :1.1 //
 
//  START 
// CELL FD3QHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD3QHSX4_SD_F_Q_R 0.1
`define FD3QHSX4_CD_F_Q_F 0.1
`define FD3QHSX4_CD_R_Q_R 0.1
`define FD3QHSX4_CP_R_Q_R 0.1
`define FD3QHSX4_CP_R_Q_F 0.1
`define FD3QHSX4_D_CP_HOLD_posedge_posedge 0.1
`define FD3QHSX4_D_CP_HOLD_negedge_posedge 0.1
`define FD3QHSX4_D_CP_SETUP_posedge_posedge 0.1
`define FD3QHSX4_D_CP_SETUP_negedge_posedge 0.1
`define FD3QHSX4_CP_PWL 0.1
`define FD3QHSX4_CP_PWH 0.1
`define FD3QHSX4_SD_PWL 0.1
`define FD3QHSX4_CD_PWL 0.1
`define FD3QHSX4_SD_CP_REC_posedge_posedge 0.1
`define FD3QHSX4_CD_CP_REC_posedge_posedge 0.1
`define FD3QHSX4_SD_CP_REM_posedge_posedge 0.1
`define FD3QHSX4_CD_CP_REM_posedge_posedge 0.1
`define FD3QHSX4_CD_SD_REC_posedge_posedge 0.1
`define FD3QHSX4_CD_SD_REM_posedge_posedge 0.1

module FD3QHSX4 (Q, D, CP, CD, SD);

   output Q;
   input D;
   input CP;
   input CD;
   input SD;


   reg Notifier;


   U_FD_P_RN_SN_NOTI u0 (IQ, D, CP, CD, SD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   and  (AndCDSD_, CD, SD);
 
   and  (AndSDD, SD, D);
   not  (D_, D);
   and  (AndCDD_, CD, D_);

   specify
`ifdef verifault

      if(CD && SD) (posedge CP => (Q +: D)) = (`FD3QHSX4_CP_R_Q_R, `FD3QHSX4_CP_R_Q_F);
      if(!SD) (posedge CD => (Q +: 1'b1)) = (`FD3QHSX4_CD_R_Q_R,`FD3QHSX4_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3QHSX4_CD_R_Q_R,`FD3QHSX4_CD_F_Q_F);
      if(CD) (negedge SD => (Q +: 1'b1)) = (`FD3QHSX4_SD_F_Q_R,`FD3QHSX4_SD_F_Q_R);

	$setuphold(posedge CP &&& AndCDSD_, posedge D, `FD3QHSX4_D_CP_SETUP_posedge_posedge, `FD3QHSX4_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSD_, negedge D, `FD3QHSX4_D_CP_SETUP_negedge_posedge, `FD3QHSX4_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD3QHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3QHSX4_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3QHSX4_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3QHSX4_CD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& AndCDD_, `FD3QHSX4_SD_CP_REC_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge CP &&& AndSDD, `FD3QHSX4_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndCDD_, posedge SD, `FD3QHSX4_SD_CP_REM_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndSDD, posedge CD, `FD3QHSX4_CD_CP_REM_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge SD, `FD3QHSX4_CD_SD_REC_posedge_posedge, Notifier);

	$hold(posedge SD, posedge CD, `FD3QHSX4_CD_SD_REM_posedge_posedge, Notifier);
`else
      (posedge CP => (Q +: D)) = (`FD3QHSX4_CP_R_Q_R, `FD3QHSX4_CP_R_Q_F);
      (posedge CD => (Q +: 1'b1)) = (`FD3QHSX4_CD_R_Q_R,`FD3QHSX4_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3QHSX4_CD_R_Q_R,`FD3QHSX4_CD_F_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD3QHSX4_SD_F_Q_R,`FD3QHSX4_SD_F_Q_R);
 
        $setuphold(posedge CP &&& AndCDSD_, posedge D, `FD3QHSX4_D_CP_SETUP_posedge_posedge, `FD3QHSX4_D_CP_HOLD_posedge_posedge, Notifier);
 $setuphold(posedge CP &&& AndCDSD_, negedge D, `FD3QHSX4_D_CP_SETUP_negedge_posedge, `FD3QHSX4_D_CP_HOLD_negedge_posedge, Notifier);
      $width(negedge CP, `FD3QHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3QHSX4_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3QHSX4_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3QHSX4_CD_PWL, 0, Notifier);
      $recovery(posedge SD, posedge CP &&& AndCDD_, `FD3QHSX4_SD_CP_REC_posedge_posedge, Notifier);
 
   $recovery(posedge CD, posedge CP &&& AndSDD, `FD3QHSX4_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndCDD_, posedge SD, `FD3QHSX4_SD_CP_REM_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndSDD, posedge CD, `FD3QHSX4_CD_CP_REM_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge SD, `FD3QHSX4_CD_SD_REC_posedge_posedge, Notifier);
 
        $hold(posedge SD, posedge CD, `FD3QHSX4_CD_SD_REM_posedge_posedge, Notifier);
 
 
`endif

   endspecify
`endif


endmodule // FD3QHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:02 and Version :1.1 //
 
//  START 
// CELL FD3SHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD3SHS_SD_F_QN_F 0.1
`define FD3SHS_CD_F_QN_R 0.1
`define FD3SHS_CD_R_QN_F 0.1
`define FD3SHS_CP_R_QN_F 0.1
`define FD3SHS_CP_R_QN_R 0.1
`define FD3SHS_SD_F_Q_R 0.1
`define FD3SHS_CD_F_Q_F 0.1
`define FD3SHS_CD_R_Q_R 0.1
`define FD3SHS_CP_R_Q_R 0.1
`define FD3SHS_CP_R_Q_F 0.1
`define FD3SHS_CD_SD_REM_posedge_posedge 0.1
`define FD3SHS_CD_SD_REC_posedge_posedge 0.1
`define FD3SHS_CD_CP_REM_posedge_posedge 0.1
`define FD3SHS_SD_CP_REM_posedge_posedge 0.1
`define FD3SHS_CD_CP_REC_posedge_posedge 0.1
`define FD3SHS_SD_CP_REC_posedge_posedge 0.1
`define FD3SHS_CD_PWL 0.1
`define FD3SHS_SD_PWL 0.1
`define FD3SHS_CP_PWH 0.1
`define FD3SHS_CP_PWL 0.1
`define FD3SHS_D_CP_SETUP_posedge_posedge 0.1
`define FD3SHS_D_CP_SETUP_negedge_posedge 0.1
`define FD3SHS_D_CP_HOLD_posedge_posedge 0.1
`define FD3SHS_D_CP_HOLD_negedge_posedge 0.1
`define FD3SHS_TI_CP_SETUP_posedge_posedge 0.1
`define FD3SHS_TI_CP_SETUP_negedge_posedge 0.1
`define FD3SHS_TI_CP_HOLD_posedge_posedge 0.1
`define FD3SHS_TI_CP_HOLD_negedge_posedge 0.1
`define FD3SHS_TE_CP_SETUP_posedge_posedge 0.1
`define FD3SHS_TE_CP_SETUP_negedge_posedge 0.1
`define FD3SHS_TE_CP_HOLD_posedge_posedge 0.1
`define FD3SHS_TE_CP_HOLD_negedge_posedge 0.1

module FD3SHS (Q, QN, D, CP, CD, SD, TI, TE);

   output Q;
   output QN;
   input D;
   input CP;
   input CD;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_SN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, SD, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   and  (AndCDSD_, CD, SD);
   and  (AndCDSDTEX_, CD, SD, TEX);
   not  (TEX, TE);
   and  (AndCDSDTE_, CD, SD, TE);
   and  (AndXorDTI_CDSD_, XorDTI_, CD, SD);
   xor  (XorDTI_, D, TI);
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);
 
   not  (D_orTI_onTE, DorTIonTE);
 
   and  (AndSDDorTI, SD, DorTIonTE);
   and  (AndCDD_orTI_, CD, D_orTI_onTE);

   specify
`ifdef verifault
      if(!TE && CD && SD) (posedge CP => (Q +: D)) = (`FD3SHS_CP_R_Q_R, `FD3SHS_CP_R_Q_F);
      if(TE && CD && SD) (posedge CP => (Q +: TI)) = (`FD3SHS_CP_R_Q_R, `FD3SHS_CP_R_Q_F);
      if(!D && TI && CD && SD) (posedge CP => (Q +: TE)) = (`FD3SHS_CP_R_Q_R, `FD3SHS_CP_R_Q_F);
      if(!TI && D && CD && SD) (posedge CP => (Q -: TE)) = (`FD3SHS_CP_R_Q_R, `FD3SHS_CP_R_Q_F);
      if(!TE && CD && SD) (posedge CP => (QN -: D)) = (`FD3SHS_CP_R_QN_R, `FD3SHS_CP_R_QN_F);
      if(TE && CD && SD) (posedge CP => (QN -: TI)) = (`FD3SHS_CP_R_QN_R, `FD3SHS_CP_R_QN_F);
      if(!D && TI && CD && SD) (posedge CP => (QN -: TE)) = (`FD3SHS_CP_R_QN_R, `FD3SHS_CP_R_QN_F);
      if(!TI && D && CD && SD) (posedge CP => (QN +: TE)) = (`FD3SHS_CP_R_QN_R, `FD3SHS_CP_R_QN_F);
      if(!SD) (posedge CD => (Q +: 1'b1)) = (`FD3SHS_CD_R_Q_R,`FD3SHS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3SHS_CD_R_Q_R,`FD3SHS_CD_F_Q_F);
      if(CD) (negedge SD => (Q +: 1'b1)) = (`FD3SHS_SD_F_Q_R,`FD3SHS_SD_F_Q_R);
      if(!SD) (posedge CD => (QN +: 1'b0)) = (`FD3SHS_CD_F_QN_R,`FD3SHS_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`FD3SHS_CD_F_QN_R,`FD3SHS_CD_R_QN_F);
      if(CD) (negedge SD => (QN +: 1'b0)) = (`FD3SHS_SD_F_QN_F,`FD3SHS_SD_F_QN_F);

	$setuphold(posedge CP &&& AndXorDTI_CDSD_, posedge TE, `FD3SHS_TE_CP_SETUP_posedge_posedge, `FD3SHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CDSD_, negedge TE, `FD3SHS_TE_CP_SETUP_negedge_posedge, `FD3SHS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDSDTE_, posedge TI, `FD3SHS_TI_CP_SETUP_posedge_posedge, `FD3SHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSDTE_, negedge TI, `FD3SHS_TI_CP_SETUP_negedge_posedge, `FD3SHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDSDTEX_, posedge D, `FD3SHS_D_CP_SETUP_posedge_posedge, `FD3SHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSDTEX_, negedge D, `FD3SHS_D_CP_SETUP_negedge_posedge, `FD3SHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD3SHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3SHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3SHS_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3SHS_CD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& AndCDD_orTI_, `FD3SHS_SD_CP_REC_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge CP &&& AndSDDorTI, `FD3SHS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndCDD_orTI_, posedge SD, `FD3SHS_SD_CP_REM_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndSDDorTI, posedge CD, `FD3SHS_CD_CP_REM_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge SD, `FD3SHS_CD_SD_REC_posedge_posedge, Notifier);

	$hold(posedge SD, posedge CD, `FD3SHS_CD_SD_REM_posedge_posedge, Notifier);
`else
       (posedge CP => (Q +: Mux21DTITE_)) = (`FD3SHS_CP_R_Q_R, `FD3SHS_CP_R_Q_F);
      (posedge CP => (QN -: Mux21DTITE_)) = (`FD3SHS_CP_R_QN_R, `FD3SHS_CP_R_QN_F);
       (posedge CD => (Q +: 1'b1)) = (`FD3SHS_CD_R_Q_R,`FD3SHS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3SHS_CD_R_Q_R,`FD3SHS_CD_F_Q_F);
       (negedge SD => (Q +: 1'b1)) = (`FD3SHS_SD_F_Q_R,`FD3SHS_SD_F_Q_R);
       (posedge CD => (QN +: 1'b0)) = (`FD3SHS_CD_F_QN_R,`FD3SHS_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`FD3SHS_CD_F_QN_R,`FD3SHS_CD_R_QN_F);
      (negedge SD => (QN +: 1'b0)) = (`FD3SHS_SD_F_QN_F,`FD3SHS_SD_F_QN_F);
 
        $setuphold(posedge CP &&& AndXorDTI_CDSD_, posedge TE, `FD3SHS_TE_CP_SETUP_posedge_posedge, `FD3SHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CDSD_, negedge TE, `FD3SHS_TE_CP_SETUP_negedge_posedge, `FD3SHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDSDTE_, posedge TI, `FD3SHS_TI_CP_SETUP_posedge_posedge, `FD3SHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSDTE_, negedge TI, `FD3SHS_TI_CP_SETUP_negedge_posedge, `FD3SHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDSDTEX_, posedge D, `FD3SHS_D_CP_SETUP_posedge_posedge, `FD3SHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSDTEX_, negedge D, `FD3SHS_D_CP_SETUP_negedge_posedge, `FD3SHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD3SHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3SHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3SHS_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3SHS_CD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& AndCDD_orTI_, `FD3SHS_SD_CP_REC_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge CP &&& AndSDDorTI, `FD3SHS_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndCDD_orTI_, posedge SD, `FD3SHS_SD_CP_REM_posedge_posedge, Notifier);
         $hold(posedge CP &&& AndSDDorTI, posedge CD, `FD3SHS_CD_CP_REM_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge SD, `FD3SHS_CD_SD_REC_posedge_posedge, Notifier);
 
        $hold(posedge SD, posedge CD, `FD3SHS_CD_SD_REM_posedge_posedge, Notifier);
 
`endif

   endspecify
`endif


endmodule // FD3SHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:04 and Version :1.1 //
 
//  START 
// CELL FD3SHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD3SHSP_SD_F_QN_F 0.1
`define FD3SHSP_CD_F_QN_R 0.1
`define FD3SHSP_CD_R_QN_F 0.1
`define FD3SHSP_CP_R_QN_F 0.1
`define FD3SHSP_CP_R_QN_R 0.1
`define FD3SHSP_SD_F_Q_R 0.1
`define FD3SHSP_CD_F_Q_F 0.1
`define FD3SHSP_CD_R_Q_R 0.1
`define FD3SHSP_CP_R_Q_R 0.1
`define FD3SHSP_CP_R_Q_F 0.1
`define FD3SHSP_CD_SD_REM_posedge_posedge 0.1
`define FD3SHSP_CD_SD_REC_posedge_posedge 0.1
`define FD3SHSP_CD_CP_REM_posedge_posedge 0.1
`define FD3SHSP_SD_CP_REM_posedge_posedge 0.1
`define FD3SHSP_CD_CP_REC_posedge_posedge 0.1
`define FD3SHSP_SD_CP_REC_posedge_posedge 0.1
`define FD3SHSP_CD_PWL 0.1
`define FD3SHSP_SD_PWL 0.1
`define FD3SHSP_CP_PWH 0.1
`define FD3SHSP_CP_PWL 0.1
`define FD3SHSP_D_CP_SETUP_posedge_posedge 0.1
`define FD3SHSP_D_CP_SETUP_negedge_posedge 0.1
`define FD3SHSP_D_CP_HOLD_posedge_posedge 0.1
`define FD3SHSP_D_CP_HOLD_negedge_posedge 0.1
`define FD3SHSP_TI_CP_SETUP_posedge_posedge 0.1
`define FD3SHSP_TI_CP_SETUP_negedge_posedge 0.1
`define FD3SHSP_TI_CP_HOLD_posedge_posedge 0.1
`define FD3SHSP_TI_CP_HOLD_negedge_posedge 0.1
`define FD3SHSP_TE_CP_SETUP_posedge_posedge 0.1
`define FD3SHSP_TE_CP_SETUP_negedge_posedge 0.1
`define FD3SHSP_TE_CP_HOLD_posedge_posedge 0.1
`define FD3SHSP_TE_CP_HOLD_negedge_posedge 0.1

module FD3SHSP (Q, QN, D, CP, CD, SD, TI, TE);

   output Q;
   output QN;
   input D;
   input CP;
   input CD;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_SN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, SD, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   and  (AndCDSD_, CD, SD);
   and  (AndCDSDTEX_, CD, SD, TEX);
   not  (TEX, TE);
   and  (AndCDSDTE_, CD, SD, TE);
   and  (AndXorDTI_CDSD_, XorDTI_, CD, SD);
   xor  (XorDTI_, D, TI);
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);
 
   not  (D_orTI_onTE, DorTIonTE);
 
   and  (AndSDDorTI, SD, DorTIonTE);
   and  (AndCDD_orTI_, CD, D_orTI_onTE);

   specify
`ifdef verifault
      if(!TE && CD && SD) (posedge CP => (Q +: D)) = (`FD3SHSP_CP_R_Q_R, `FD3SHSP_CP_R_Q_F);
      if(TE && CD && SD) (posedge CP => (Q +: TI)) = (`FD3SHSP_CP_R_Q_R, `FD3SHSP_CP_R_Q_F);
      if(!D && TI && CD && SD) (posedge CP => (Q +: TE)) = (`FD3SHSP_CP_R_Q_R, `FD3SHSP_CP_R_Q_F);
      if(!TI && D && CD && SD) (posedge CP => (Q -: TE)) = (`FD3SHSP_CP_R_Q_R, `FD3SHSP_CP_R_Q_F);
      if(!TE && CD && SD) (posedge CP => (QN -: D)) = (`FD3SHSP_CP_R_QN_R, `FD3SHSP_CP_R_QN_F);
      if(TE && CD && SD) (posedge CP => (QN -: TI)) = (`FD3SHSP_CP_R_QN_R, `FD3SHSP_CP_R_QN_F);
      if(!D && TI && CD && SD) (posedge CP => (QN -: TE)) = (`FD3SHSP_CP_R_QN_R, `FD3SHSP_CP_R_QN_F);
      if(!TI && D && CD && SD) (posedge CP => (QN +: TE)) = (`FD3SHSP_CP_R_QN_R, `FD3SHSP_CP_R_QN_F);
      if(!SD) (posedge CD => (Q +: 1'b1)) = (`FD3SHSP_CD_R_Q_R,`FD3SHSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3SHSP_CD_R_Q_R,`FD3SHSP_CD_F_Q_F);
      if(CD) (negedge SD => (Q +: 1'b1)) = (`FD3SHSP_SD_F_Q_R,`FD3SHSP_SD_F_Q_R);
      if(!SD) (posedge CD => (QN +: 1'b0)) = (`FD3SHSP_CD_F_QN_R,`FD3SHSP_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`FD3SHSP_CD_F_QN_R,`FD3SHSP_CD_R_QN_F);
      if(CD) (negedge SD => (QN +: 1'b0)) = (`FD3SHSP_SD_F_QN_F,`FD3SHSP_SD_F_QN_F);

	$setuphold(posedge CP &&& AndXorDTI_CDSD_, posedge TE, `FD3SHSP_TE_CP_SETUP_posedge_posedge, `FD3SHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CDSD_, negedge TE, `FD3SHSP_TE_CP_SETUP_negedge_posedge, `FD3SHSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDSDTE_, posedge TI, `FD3SHSP_TI_CP_SETUP_posedge_posedge, `FD3SHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSDTE_, negedge TI, `FD3SHSP_TI_CP_SETUP_negedge_posedge, `FD3SHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDSDTEX_, posedge D, `FD3SHSP_D_CP_SETUP_posedge_posedge, `FD3SHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSDTEX_, negedge D, `FD3SHSP_D_CP_SETUP_negedge_posedge, `FD3SHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD3SHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3SHSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3SHSP_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3SHSP_CD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& AndCDD_orTI_, `FD3SHSP_SD_CP_REC_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge CP &&& AndSDDorTI, `FD3SHSP_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndCDD_orTI_, posedge SD, `FD3SHSP_SD_CP_REM_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndSDDorTI, posedge CD, `FD3SHSP_CD_CP_REM_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge SD, `FD3SHSP_CD_SD_REC_posedge_posedge, Notifier);

	$hold(posedge SD, posedge CD, `FD3SHSP_CD_SD_REM_posedge_posedge, Notifier);
`else
       (posedge CP => (Q +: Mux21DTITE_)) = (`FD3SHSP_CP_R_Q_R, `FD3SHSP_CP_R_Q_F);
      (posedge CP => (QN -: Mux21DTITE_)) = (`FD3SHSP_CP_R_QN_R, `FD3SHSP_CP_R_QN_F);
       (posedge CD => (Q +: 1'b1)) = (`FD3SHSP_CD_R_Q_R,`FD3SHSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3SHSP_CD_R_Q_R,`FD3SHSP_CD_F_Q_F);
       (negedge SD => (Q +: 1'b1)) = (`FD3SHSP_SD_F_Q_R,`FD3SHSP_SD_F_Q_R);
       (posedge CD => (QN +: 1'b0)) = (`FD3SHSP_CD_F_QN_R,`FD3SHSP_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`FD3SHSP_CD_F_QN_R,`FD3SHSP_CD_R_QN_F);
      (negedge SD => (QN +: 1'b0)) = (`FD3SHSP_SD_F_QN_F,`FD3SHSP_SD_F_QN_F);
 
        $setuphold(posedge CP &&& AndXorDTI_CDSD_, posedge TE, `FD3SHSP_TE_CP_SETUP_posedge_posedge, `FD3SHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CDSD_, negedge TE, `FD3SHSP_TE_CP_SETUP_negedge_posedge, `FD3SHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDSDTE_, posedge TI, `FD3SHSP_TI_CP_SETUP_posedge_posedge, `FD3SHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSDTE_, negedge TI, `FD3SHSP_TI_CP_SETUP_negedge_posedge, `FD3SHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDSDTEX_, posedge D, `FD3SHSP_D_CP_SETUP_posedge_posedge, `FD3SHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSDTEX_, negedge D, `FD3SHSP_D_CP_SETUP_negedge_posedge, `FD3SHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD3SHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3SHSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3SHSP_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3SHSP_CD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& AndCDD_orTI_, `FD3SHSP_SD_CP_REC_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge CP &&& AndSDDorTI, `FD3SHSP_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndCDD_orTI_, posedge SD, `FD3SHSP_SD_CP_REM_posedge_posedge, Notifier);
         $hold(posedge CP &&& AndSDDorTI, posedge CD, `FD3SHSP_CD_CP_REM_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge SD, `FD3SHSP_CD_SD_REC_posedge_posedge, Notifier);
 
        $hold(posedge SD, posedge CD, `FD3SHSP_CD_SD_REM_posedge_posedge, Notifier);
 
`endif

   endspecify
`endif


endmodule // FD3SHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:04 and Version :1.1 //
 
//  START 
// CELL FD3SQHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD3SQHS_SD_F_Q_R 0.1
`define FD3SQHS_CD_F_Q_F 0.1
`define FD3SQHS_CD_R_Q_R 0.1
`define FD3SQHS_CP_R_Q_R 0.1
`define FD3SQHS_CP_R_Q_F 0.1
`define FD3SQHS_TE_CP_HOLD_posedge_posedge 0.1
`define FD3SQHS_TE_CP_HOLD_negedge_posedge 0.1
`define FD3SQHS_TE_CP_SETUP_posedge_posedge 0.1
`define FD3SQHS_TE_CP_SETUP_negedge_posedge 0.1
`define FD3SQHS_TI_CP_HOLD_posedge_posedge 0.1
`define FD3SQHS_TI_CP_HOLD_negedge_posedge 0.1
`define FD3SQHS_TI_CP_SETUP_posedge_posedge 0.1
`define FD3SQHS_TI_CP_SETUP_negedge_posedge 0.1
`define FD3SQHS_D_CP_HOLD_posedge_posedge 0.1
`define FD3SQHS_D_CP_HOLD_negedge_posedge 0.1
`define FD3SQHS_D_CP_SETUP_posedge_posedge 0.1
`define FD3SQHS_D_CP_SETUP_negedge_posedge 0.1
`define FD3SQHS_CP_PWL 0.1
`define FD3SQHS_CP_PWH 0.1
`define FD3SQHS_SD_PWL 0.1
`define FD3SQHS_CD_PWL 0.1
`define FD3SQHS_SD_CP_REC_posedge_posedge 0.1
`define FD3SQHS_CD_CP_REC_posedge_posedge 0.1
`define FD3SQHS_SD_CP_REM_posedge_posedge 0.1
`define FD3SQHS_CD_CP_REM_posedge_posedge 0.1
`define FD3SQHS_CD_SD_REC_posedge_posedge 0.1
`define FD3SQHS_CD_SD_REM_posedge_posedge 0.1

module FD3SQHS (Q, D, CP, CD, SD, TI, TE);

   output Q;
   input D;
   input CP;
   input CD;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_SN_NOTI u1 (IQ, Mux21DTITE_, CP, CD, SD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   and  (AndCDSD_, CD, SD);
   and  (AndCDSDTEX_, CD, SD, TEX);
   not  (TEX, TE);
   and  (AndCDSDTE_, CD, SD, TE);
   and  (AndXorDTI_CDSD_, XorDTI_, CD, SD);
   xor  (XorDTI_, D, TI);
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);
 
   not  (D_orTI_onTE, DorTIonTE);
 
   and  (AndSDDorTI, SD, DorTIonTE);
   and  (AndCDD_orTI_, CD, D_orTI_onTE);

   specify
`ifdef verifault 
      if(!TE && CD && SD) (posedge CP => (Q +: D)) = (`FD3SQHS_CP_R_Q_R, `FD3SQHS_CP_R_Q_F);
      if(TE && CD && SD) (posedge CP => (Q +: TI)) = (`FD3SQHS_CP_R_Q_R, `FD3SQHS_CP_R_Q_F);
      if(!D && TI && CD && SD) (posedge CP => (Q +: TE)) = (`FD3SQHS_CP_R_Q_R, `FD3SQHS_CP_R_Q_F);
      if(!TI && D && CD && SD) (posedge CP => (Q -: TE)) = (`FD3SQHS_CP_R_Q_R, `FD3SQHS_CP_R_Q_F);
      if(!SD) (posedge CD => (Q +: 1'b1)) = (`FD3SQHS_CD_R_Q_R,`FD3SQHS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3SQHS_CD_R_Q_R,`FD3SQHS_CD_F_Q_F);
      if(CD) (negedge SD => (Q +: 1'b1)) = (`FD3SQHS_SD_F_Q_R,`FD3SQHS_SD_F_Q_R);

	$setuphold(posedge CP &&& AndXorDTI_CDSD_, posedge TE, `FD3SQHS_TE_CP_SETUP_posedge_posedge, `FD3SQHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CDSD_, negedge TE, `FD3SQHS_TE_CP_SETUP_negedge_posedge, `FD3SQHS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDSDTE_, posedge TI, `FD3SQHS_TI_CP_SETUP_posedge_posedge, `FD3SQHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSDTE_, negedge TI, `FD3SQHS_TI_CP_SETUP_negedge_posedge, `FD3SQHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDSDTEX_, posedge D, `FD3SQHS_D_CP_SETUP_posedge_posedge, `FD3SQHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSDTEX_, negedge D, `FD3SQHS_D_CP_SETUP_negedge_posedge, `FD3SQHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD3SQHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3SQHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3SQHS_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3SQHS_CD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& AndCDD_orTI_, `FD3SQHS_SD_CP_REC_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge CP &&& AndSDDorTI, `FD3SQHS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndCDD_orTI_, posedge SD, `FD3SQHS_SD_CP_REM_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndSDDorTI, posedge CD, `FD3SQHS_CD_CP_REM_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge SD, `FD3SQHS_CD_SD_REC_posedge_posedge, Notifier);

	$hold(posedge SD, posedge CD, `FD3SQHS_CD_SD_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FD3SQHS_CP_R_Q_R, `FD3SQHS_CP_R_Q_F);
      (posedge CD => (Q +: 1'b1)) = (`FD3SQHS_CD_R_Q_R,`FD3SQHS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3SQHS_CD_R_Q_R,`FD3SQHS_CD_F_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD3SQHS_SD_F_Q_R,`FD3SQHS_SD_F_Q_R);
 
        $setuphold(posedge CP &&& AndXorDTI_CDSD_, posedge TE, `FD3SQHS_TE_CP_SETUP_posedge_posedge, `FD3SQHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CDSD_, negedge TE, `FD3SQHS_TE_CP_SETUP_negedge_posedge, `FD3SQHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDSDTE_, posedge TI, `FD3SQHS_TI_CP_SETUP_posedge_posedge, `FD3SQHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSDTE_, negedge TI, `FD3SQHS_TI_CP_SETUP_negedge_posedge, `FD3SQHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDSDTEX_, posedge D, `FD3SQHS_D_CP_SETUP_posedge_posedge, `FD3SQHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSDTEX_, negedge D, `FD3SQHS_D_CP_SETUP_negedge_posedge, `FD3SQHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD3SQHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3SQHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3SQHS_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3SQHS_CD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& AndCDD_orTI_, `FD3SQHS_SD_CP_REC_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge CP &&& AndSDDorTI, `FD3SQHS_CD_CP_REC_posedge_posedge,Notifier);
 
        $hold(posedge CP &&& AndCDD_orTI_, posedge SD, `FD3SQHS_SD_CP_REM_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndSDDorTI, posedge CD, `FD3SQHS_CD_CP_REM_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge SD, `FD3SQHS_CD_SD_REC_posedge_posedge, Notifier);
 
        $hold(posedge SD, posedge CD, `FD3SQHS_CD_SD_REM_posedge_posedge, Notifier);
 
 
`endif
   endspecify
`endif


endmodule // FD3SQHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:08 and Version :1.1 //
 
//  START 
// CELL FD3SQHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD3SQHSP_SD_F_Q_R 0.1
`define FD3SQHSP_CD_F_Q_F 0.1
`define FD3SQHSP_CD_R_Q_R 0.1
`define FD3SQHSP_CP_R_Q_R 0.1
`define FD3SQHSP_CP_R_Q_F 0.1
`define FD3SQHSP_TE_CP_HOLD_posedge_posedge 0.1
`define FD3SQHSP_TE_CP_HOLD_negedge_posedge 0.1
`define FD3SQHSP_TE_CP_SETUP_posedge_posedge 0.1
`define FD3SQHSP_TE_CP_SETUP_negedge_posedge 0.1
`define FD3SQHSP_TI_CP_HOLD_posedge_posedge 0.1
`define FD3SQHSP_TI_CP_HOLD_negedge_posedge 0.1
`define FD3SQHSP_TI_CP_SETUP_posedge_posedge 0.1
`define FD3SQHSP_TI_CP_SETUP_negedge_posedge 0.1
`define FD3SQHSP_D_CP_HOLD_posedge_posedge 0.1
`define FD3SQHSP_D_CP_HOLD_negedge_posedge 0.1
`define FD3SQHSP_D_CP_SETUP_posedge_posedge 0.1
`define FD3SQHSP_D_CP_SETUP_negedge_posedge 0.1
`define FD3SQHSP_CP_PWL 0.1
`define FD3SQHSP_CP_PWH 0.1
`define FD3SQHSP_SD_PWL 0.1
`define FD3SQHSP_CD_PWL 0.1
`define FD3SQHSP_SD_CP_REC_posedge_posedge 0.1
`define FD3SQHSP_CD_CP_REC_posedge_posedge 0.1
`define FD3SQHSP_SD_CP_REM_posedge_posedge 0.1
`define FD3SQHSP_CD_CP_REM_posedge_posedge 0.1
`define FD3SQHSP_CD_SD_REC_posedge_posedge 0.1
`define FD3SQHSP_CD_SD_REM_posedge_posedge 0.1

module FD3SQHSP (Q, D, CP, CD, SD, TI, TE);

   output Q;
   input D;
   input CP;
   input CD;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_SN_NOTI u1 (IQ, Mux21DTITE_, CP, CD, SD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   and  (AndCDSD_, CD, SD);
   and  (AndCDSDTEX_, CD, SD, TEX);
   not  (TEX, TE);
   and  (AndCDSDTE_, CD, SD, TE);
   and  (AndXorDTI_CDSD_, XorDTI_, CD, SD);
   xor  (XorDTI_, D, TI);
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);
 
   not  (D_orTI_onTE, DorTIonTE);
 
   and  (AndSDDorTI, SD, DorTIonTE);
   and  (AndCDD_orTI_, CD, D_orTI_onTE);

   specify
`ifdef verifault 
      if(!TE && CD && SD) (posedge CP => (Q +: D)) = (`FD3SQHSP_CP_R_Q_R, `FD3SQHSP_CP_R_Q_F);
      if(TE && CD && SD) (posedge CP => (Q +: TI)) = (`FD3SQHSP_CP_R_Q_R, `FD3SQHSP_CP_R_Q_F);
      if(!D && TI && CD && SD) (posedge CP => (Q +: TE)) = (`FD3SQHSP_CP_R_Q_R, `FD3SQHSP_CP_R_Q_F);
      if(!TI && D && CD && SD) (posedge CP => (Q -: TE)) = (`FD3SQHSP_CP_R_Q_R, `FD3SQHSP_CP_R_Q_F);
      if(!SD) (posedge CD => (Q +: 1'b1)) = (`FD3SQHSP_CD_R_Q_R,`FD3SQHSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3SQHSP_CD_R_Q_R,`FD3SQHSP_CD_F_Q_F);
      if(CD) (negedge SD => (Q +: 1'b1)) = (`FD3SQHSP_SD_F_Q_R,`FD3SQHSP_SD_F_Q_R);

	$setuphold(posedge CP &&& AndXorDTI_CDSD_, posedge TE, `FD3SQHSP_TE_CP_SETUP_posedge_posedge, `FD3SQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CDSD_, negedge TE, `FD3SQHSP_TE_CP_SETUP_negedge_posedge, `FD3SQHSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDSDTE_, posedge TI, `FD3SQHSP_TI_CP_SETUP_posedge_posedge, `FD3SQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSDTE_, negedge TI, `FD3SQHSP_TI_CP_SETUP_negedge_posedge, `FD3SQHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDSDTEX_, posedge D, `FD3SQHSP_D_CP_SETUP_posedge_posedge, `FD3SQHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSDTEX_, negedge D, `FD3SQHSP_D_CP_SETUP_negedge_posedge, `FD3SQHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD3SQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3SQHSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3SQHSP_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3SQHSP_CD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& AndCDD_orTI_, `FD3SQHSP_SD_CP_REC_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge CP &&& AndSDDorTI, `FD3SQHSP_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndCDD_orTI_, posedge SD, `FD3SQHSP_SD_CP_REM_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndSDDorTI, posedge CD, `FD3SQHSP_CD_CP_REM_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge SD, `FD3SQHSP_CD_SD_REC_posedge_posedge, Notifier);

	$hold(posedge SD, posedge CD, `FD3SQHSP_CD_SD_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FD3SQHSP_CP_R_Q_R, `FD3SQHSP_CP_R_Q_F);
      (posedge CD => (Q +: 1'b1)) = (`FD3SQHSP_CD_R_Q_R,`FD3SQHSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3SQHSP_CD_R_Q_R,`FD3SQHSP_CD_F_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD3SQHSP_SD_F_Q_R,`FD3SQHSP_SD_F_Q_R);
 
        $setuphold(posedge CP &&& AndXorDTI_CDSD_, posedge TE, `FD3SQHSP_TE_CP_SETUP_posedge_posedge, `FD3SQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CDSD_, negedge TE, `FD3SQHSP_TE_CP_SETUP_negedge_posedge, `FD3SQHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDSDTE_, posedge TI, `FD3SQHSP_TI_CP_SETUP_posedge_posedge, `FD3SQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSDTE_, negedge TI, `FD3SQHSP_TI_CP_SETUP_negedge_posedge, `FD3SQHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDSDTEX_, posedge D, `FD3SQHSP_D_CP_SETUP_posedge_posedge, `FD3SQHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSDTEX_, negedge D, `FD3SQHSP_D_CP_SETUP_negedge_posedge, `FD3SQHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD3SQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3SQHSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3SQHSP_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3SQHSP_CD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& AndCDD_orTI_, `FD3SQHSP_SD_CP_REC_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge CP &&& AndSDDorTI, `FD3SQHSP_CD_CP_REC_posedge_posedge,Notifier);
 
        $hold(posedge CP &&& AndCDD_orTI_, posedge SD, `FD3SQHSP_SD_CP_REM_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndSDDorTI, posedge CD, `FD3SQHSP_CD_CP_REM_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge SD, `FD3SQHSP_CD_SD_REC_posedge_posedge, Notifier);
 
        $hold(posedge SD, posedge CD, `FD3SQHSP_CD_SD_REM_posedge_posedge, Notifier);
 
 
`endif
   endspecify
`endif


endmodule // FD3SQHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:08 and Version :1.1 //
 
//  START 
// CELL FD3SQHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD3SQHSX4_SD_F_Q_R 0.1
`define FD3SQHSX4_CD_F_Q_F 0.1
`define FD3SQHSX4_CD_R_Q_R 0.1
`define FD3SQHSX4_CP_R_Q_R 0.1
`define FD3SQHSX4_CP_R_Q_F 0.1
`define FD3SQHSX4_TE_CP_HOLD_posedge_posedge 0.1
`define FD3SQHSX4_TE_CP_HOLD_negedge_posedge 0.1
`define FD3SQHSX4_TE_CP_SETUP_posedge_posedge 0.1
`define FD3SQHSX4_TE_CP_SETUP_negedge_posedge 0.1
`define FD3SQHSX4_TI_CP_HOLD_posedge_posedge 0.1
`define FD3SQHSX4_TI_CP_HOLD_negedge_posedge 0.1
`define FD3SQHSX4_TI_CP_SETUP_posedge_posedge 0.1
`define FD3SQHSX4_TI_CP_SETUP_negedge_posedge 0.1
`define FD3SQHSX4_D_CP_HOLD_posedge_posedge 0.1
`define FD3SQHSX4_D_CP_HOLD_negedge_posedge 0.1
`define FD3SQHSX4_D_CP_SETUP_posedge_posedge 0.1
`define FD3SQHSX4_D_CP_SETUP_negedge_posedge 0.1
`define FD3SQHSX4_CP_PWL 0.1
`define FD3SQHSX4_CP_PWH 0.1
`define FD3SQHSX4_SD_PWL 0.1
`define FD3SQHSX4_CD_PWL 0.1
`define FD3SQHSX4_SD_CP_REC_posedge_posedge 0.1
`define FD3SQHSX4_CD_CP_REC_posedge_posedge 0.1
`define FD3SQHSX4_SD_CP_REM_posedge_posedge 0.1
`define FD3SQHSX4_CD_CP_REM_posedge_posedge 0.1
`define FD3SQHSX4_CD_SD_REC_posedge_posedge 0.1
`define FD3SQHSX4_CD_SD_REM_posedge_posedge 0.1

module FD3SQHSX4 (Q, D, CP, CD, SD, TI, TE);

   output Q;
   input D;
   input CP;
   input CD;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_SN_NOTI u1 (IQ, Mux21DTITE_, CP, CD, SD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   and  (AndCDSD_, CD, SD);
   and  (AndCDSDTEX_, CD, SD, TEX);
   not  (TEX, TE);
   and  (AndCDSDTE_, CD, SD, TE);
   and  (AndXorDTI_CDSD_, XorDTI_, CD, SD);
   xor  (XorDTI_, D, TI);
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);
 
   not  (D_orTI_onTE, DorTIonTE);
 
   and  (AndSDDorTI, SD, DorTIonTE);
   and  (AndCDD_orTI_, CD, D_orTI_onTE);

   specify
`ifdef verifault 
      if(!TE && CD && SD) (posedge CP => (Q +: D)) = (`FD3SQHSX4_CP_R_Q_R, `FD3SQHSX4_CP_R_Q_F);
      if(TE && CD && SD) (posedge CP => (Q +: TI)) = (`FD3SQHSX4_CP_R_Q_R, `FD3SQHSX4_CP_R_Q_F);
      if(!D && TI && CD && SD) (posedge CP => (Q +: TE)) = (`FD3SQHSX4_CP_R_Q_R, `FD3SQHSX4_CP_R_Q_F);
      if(!TI && D && CD && SD) (posedge CP => (Q -: TE)) = (`FD3SQHSX4_CP_R_Q_R, `FD3SQHSX4_CP_R_Q_F);
      if(!SD) (posedge CD => (Q +: 1'b1)) = (`FD3SQHSX4_CD_R_Q_R,`FD3SQHSX4_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3SQHSX4_CD_R_Q_R,`FD3SQHSX4_CD_F_Q_F);
      if(CD) (negedge SD => (Q +: 1'b1)) = (`FD3SQHSX4_SD_F_Q_R,`FD3SQHSX4_SD_F_Q_R);

	$setuphold(posedge CP &&& AndXorDTI_CDSD_, posedge TE, `FD3SQHSX4_TE_CP_SETUP_posedge_posedge, `FD3SQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CDSD_, negedge TE, `FD3SQHSX4_TE_CP_SETUP_negedge_posedge, `FD3SQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDSDTE_, posedge TI, `FD3SQHSX4_TI_CP_SETUP_posedge_posedge, `FD3SQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSDTE_, negedge TI, `FD3SQHSX4_TI_CP_SETUP_negedge_posedge, `FD3SQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDSDTEX_, posedge D, `FD3SQHSX4_D_CP_SETUP_posedge_posedge, `FD3SQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSDTEX_, negedge D, `FD3SQHSX4_D_CP_SETUP_negedge_posedge, `FD3SQHSX4_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD3SQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3SQHSX4_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3SQHSX4_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3SQHSX4_CD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& AndCDD_orTI_, `FD3SQHSX4_SD_CP_REC_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge CP &&& AndSDDorTI, `FD3SQHSX4_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndCDD_orTI_, posedge SD, `FD3SQHSX4_SD_CP_REM_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndSDDorTI, posedge CD, `FD3SQHSX4_CD_CP_REM_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge SD, `FD3SQHSX4_CD_SD_REC_posedge_posedge, Notifier);

	$hold(posedge SD, posedge CD, `FD3SQHSX4_CD_SD_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FD3SQHSX4_CP_R_Q_R, `FD3SQHSX4_CP_R_Q_F);
      (posedge CD => (Q +: 1'b1)) = (`FD3SQHSX4_CD_R_Q_R,`FD3SQHSX4_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3SQHSX4_CD_R_Q_R,`FD3SQHSX4_CD_F_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD3SQHSX4_SD_F_Q_R,`FD3SQHSX4_SD_F_Q_R);
 
        $setuphold(posedge CP &&& AndXorDTI_CDSD_, posedge TE, `FD3SQHSX4_TE_CP_SETUP_posedge_posedge, `FD3SQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CDSD_, negedge TE, `FD3SQHSX4_TE_CP_SETUP_negedge_posedge, `FD3SQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDSDTE_, posedge TI, `FD3SQHSX4_TI_CP_SETUP_posedge_posedge, `FD3SQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSDTE_, negedge TI, `FD3SQHSX4_TI_CP_SETUP_negedge_posedge, `FD3SQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDSDTEX_, posedge D, `FD3SQHSX4_D_CP_SETUP_posedge_posedge, `FD3SQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSDTEX_, negedge D, `FD3SQHSX4_D_CP_SETUP_negedge_posedge, `FD3SQHSX4_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD3SQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3SQHSX4_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3SQHSX4_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3SQHSX4_CD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& AndCDD_orTI_, `FD3SQHSX4_SD_CP_REC_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge CP &&& AndSDDorTI, `FD3SQHSX4_CD_CP_REC_posedge_posedge,Notifier);
 
        $hold(posedge CP &&& AndCDD_orTI_, posedge SD, `FD3SQHSX4_SD_CP_REM_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndSDDorTI, posedge CD, `FD3SQHSX4_CD_CP_REM_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge SD, `FD3SQHSX4_CD_SD_REC_posedge_posedge, Notifier);
 
        $hold(posedge SD, posedge CD, `FD3SQHSX4_CD_SD_REM_posedge_posedge, Notifier);
 
 
`endif
   endspecify
`endif


endmodule // FD3SQHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:08 and Version :1.1 //
 
//  START 
// CELL FD3THS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD3THS_SD_F_SO_R 0.1
`define FD3THS_CD_F_SO_F 0.1
`define FD3THS_CD_R_SO_R 0.1
`define FD3THS_CP_R_SO_R 0.1
`define FD3THS_CP_R_SO_F 0.1
`define FD3THS_SD_F_QN_F 0.1
`define FD3THS_CD_F_QN_R 0.1
`define FD3THS_CD_R_QN_F 0.1
`define FD3THS_CP_R_QN_F 0.1
`define FD3THS_CP_R_QN_R 0.1
`define FD3THS_SD_F_Q_R 0.1
`define FD3THS_CD_F_Q_F 0.1
`define FD3THS_CD_R_Q_R 0.1
`define FD3THS_CP_R_Q_R 0.1
`define FD3THS_CP_R_Q_F 0.1
`define FD3THS_CD_SD_REM_posedge_posedge 0.1
`define FD3THS_CD_SD_REC_posedge_posedge 0.1
`define FD3THS_CD_CP_REM_posedge_posedge 0.1
`define FD3THS_SD_CP_REM_posedge_posedge 0.1
`define FD3THS_CD_CP_REC_posedge_posedge 0.1
`define FD3THS_SD_CP_REC_posedge_posedge 0.1
`define FD3THS_CD_PWL 0.1
`define FD3THS_SD_PWL 0.1
`define FD3THS_CP_PWH 0.1
`define FD3THS_CP_PWL 0.1
`define FD3THS_D_CP_SETUP_posedge_posedge 0.1
`define FD3THS_D_CP_SETUP_negedge_posedge 0.1
`define FD3THS_D_CP_HOLD_posedge_posedge 0.1
`define FD3THS_D_CP_HOLD_negedge_posedge 0.1
`define FD3THS_TI_CP_SETUP_posedge_posedge 0.1
`define FD3THS_TI_CP_SETUP_negedge_posedge 0.1
`define FD3THS_TI_CP_HOLD_posedge_posedge 0.1
`define FD3THS_TI_CP_HOLD_negedge_posedge 0.1
`define FD3THS_TE_CP_SETUP_posedge_posedge 0.1
`define FD3THS_TE_CP_SETUP_negedge_posedge 0.1
`define FD3THS_TE_CP_HOLD_posedge_posedge 0.1
`define FD3THS_TE_CP_HOLD_negedge_posedge 0.1

module FD3THS (Q, QN, SO, D, CP, CD, SD, TI, TE);

   output Q;
   output QN;
   output SO;
   input D;
   input CP;
   input CD;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_SN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, SD, Notifier);

   buf  u2 (Q, IQ);
   buf  u3 (SO, IQ);
   not  u4 (QN, IQ);



`ifdef functional
`else
   and  (AndCDSD_, CD, SD);
   not  (TEX, TE);
   and  (AndCDSDTEX_, CD, SD, TEX);
   and  (AndCDSDTE_, CD, SD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_CDSD_, XorDTI_, CD, SD);
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);
 
   not  (D_orTI_onTE, DorTIonTE);
 
   and  (AndSDDorTI, SD, DorTIonTE);
   and  (AndCDD_orTI_, CD, D_orTI_onTE);

   specify
`ifdef verifault

      if(!TE && CD && SD) (posedge CP => (Q +: D)) = (`FD3THS_CP_R_Q_R, `FD3THS_CP_R_Q_F);
      if(TE && CD && SD) (posedge CP => (Q +: TI)) = (`FD3THS_CP_R_Q_R, `FD3THS_CP_R_Q_F);
      if(!D && TI && CD && SD) (posedge CP => (Q +: TE)) = (`FD3THS_CP_R_Q_R, `FD3THS_CP_R_Q_F);
      if(!TI && D && CD && SD) (posedge CP => (Q -: TE)) = (`FD3THS_CP_R_Q_R, `FD3THS_CP_R_Q_F);
      if(!TE && CD && SD) (posedge CP => (QN -: D)) = (`FD3THS_CP_R_QN_R, `FD3THS_CP_R_QN_F);
      if(TE && CD && SD) (posedge CP => (QN -: TI)) = (`FD3THS_CP_R_QN_R, `FD3THS_CP_R_QN_F);
      if(!D && TI && CD && SD) (posedge CP => (QN -: TE)) = (`FD3THS_CP_R_QN_R, `FD3THS_CP_R_QN_F);
      if(!TI && D && CD && SD) (posedge CP => (QN +: TE)) = (`FD3THS_CP_R_QN_R, `FD3THS_CP_R_QN_F);
      if(!TE && CD && SD) (posedge CP => (SO +: D)) = (`FD3THS_CP_R_SO_R, `FD3THS_CP_R_SO_F);
      if(TE && CD && SD) (posedge CP => (SO +: TI)) = (`FD3THS_CP_R_SO_R, `FD3THS_CP_R_SO_F);
      if(!D && TI && CD && SD) (posedge CP => (SO +: TE)) = (`FD3THS_CP_R_SO_R, `FD3THS_CP_R_SO_F);
      if(!TI && D && CD && SD) (posedge CP => (SO -: TE)) = (`FD3THS_CP_R_SO_R, `FD3THS_CP_R_SO_F);
      if(!SD) (posedge CD => (Q +: 1'b1)) = (`FD3THS_CD_R_Q_R,`FD3THS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3THS_CD_R_Q_R,`FD3THS_CD_F_Q_F);
      if(CD) (negedge SD => (Q +: 1'b1)) = (`FD3THS_SD_F_Q_R,`FD3THS_SD_F_Q_R);
      if(!SD) (posedge CD => (QN +: 1'b0)) = (`FD3THS_CD_F_QN_R,`FD3THS_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`FD3THS_CD_F_QN_R,`FD3THS_CD_R_QN_F);
      if(CD) (negedge SD => (QN +: 1'b0)) = (`FD3THS_SD_F_QN_F,`FD3THS_SD_F_QN_F);
      if(!SD) (posedge CD => (SO +: 1'b1)) = (`FD3THS_CD_R_SO_R,`FD3THS_CD_F_SO_F);
      (negedge CD => (SO +: 1'b0)) = (`FD3THS_CD_R_SO_R,`FD3THS_CD_F_SO_F);
      if(CD) (negedge SD => (SO +: 1'b1)) = (`FD3THS_SD_F_SO_R,`FD3THS_SD_F_SO_R);

	$setuphold(posedge CP &&& AndXorDTI_CDSD_, posedge TE, `FD3THS_TE_CP_SETUP_posedge_posedge, `FD3THS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CDSD_, negedge TE, `FD3THS_TE_CP_SETUP_negedge_posedge, `FD3THS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDSDTE_, posedge TI, `FD3THS_TI_CP_SETUP_posedge_posedge, `FD3THS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSDTE_, negedge TI, `FD3THS_TI_CP_SETUP_negedge_posedge, `FD3THS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDSDTEX_, posedge D, `FD3THS_D_CP_SETUP_posedge_posedge, `FD3THS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSDTEX_, negedge D, `FD3THS_D_CP_SETUP_negedge_posedge, `FD3THS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD3THS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3THS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3THS_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3THS_CD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& AndCDD_orTI_, `FD3THS_SD_CP_REC_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge CP &&& AndSDDorTI, `FD3THS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndCDD_orTI_, posedge SD, `FD3THS_SD_CP_REM_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndSDDorTI, posedge CD, `FD3THS_CD_CP_REM_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge SD, `FD3THS_CD_SD_REC_posedge_posedge, Notifier);

	$hold(posedge SD, posedge CD, `FD3THS_CD_SD_REM_posedge_posedge, Notifier);
`else

      (posedge CP => (Q +: Mux21DTITE_)) = (`FD3THS_CP_R_Q_R, `FD3THS_CP_R_Q_F);
      (posedge CP => (QN -: Mux21DTITE_)) = (`FD3THS_CP_R_QN_R, `FD3THS_CP_R_QN_F);
      (posedge CP => (SO +: Mux21DTITE_)) = (`FD3THS_CP_R_SO_R, `FD3THS_CP_R_SO_F);
      (posedge CD => (Q +: 1'b1)) = (`FD3THS_CD_R_Q_R,`FD3THS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3THS_CD_R_Q_R,`FD3THS_CD_F_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD3THS_SD_F_Q_R,`FD3THS_SD_F_Q_R);
      (posedge CD => (QN +: 1'b0)) = (`FD3THS_CD_F_QN_R,`FD3THS_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`FD3THS_CD_F_QN_R,`FD3THS_CD_R_QN_F);
      (negedge SD => (QN +: 1'b0)) = (`FD3THS_SD_F_QN_F,`FD3THS_SD_F_QN_F);
      (posedge CD => (SO +: 1'b1)) = (`FD3THS_CD_R_SO_R,`FD3THS_CD_F_SO_F);
      (negedge CD => (SO +: 1'b0)) = (`FD3THS_CD_R_SO_R,`FD3THS_CD_F_SO_F);
      (negedge SD => (SO +: 1'b1)) = (`FD3THS_SD_F_SO_R,`FD3THS_SD_F_SO_R);
 
        $setuphold(posedge CP &&& AndXorDTI_CDSD_, posedge TE, `FD3THS_TE_CP_SETUP_posedge_posedge, `FD3THS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CDSD_, negedge TE, `FD3THS_TE_CP_SETUP_negedge_posedge, `FD3THS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDSDTE_, posedge TI, `FD3THS_TI_CP_SETUP_posedge_posedge, `FD3THS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSDTE_, negedge TI, `FD3THS_TI_CP_SETUP_negedge_posedge, `FD3THS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDSDTEX_, posedge D, `FD3THS_D_CP_SETUP_posedge_posedge, `FD3THS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSDTEX_, negedge D, `FD3THS_D_CP_SETUP_negedge_posedge, `FD3THS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD3THS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3THS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3THS_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3THS_CD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& AndCDD_orTI_, `FD3THS_SD_CP_REC_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge CP &&& AndSDDorTI, `FD3THS_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndCDD_orTI_, posedge SD, `FD3THS_SD_CP_REM_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndSDDorTI, posedge CD, `FD3THS_CD_CP_REM_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge SD, `FD3THS_CD_SD_REC_posedge_posedge, Notifier);
 
        $hold(posedge SD, posedge CD, `FD3THS_CD_SD_REM_posedge_posedge, Notifier);
`endif

   endspecify
`endif


endmodule // FD3THS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:11 and Version :1.1 //
 
//  START 
// CELL FD3THSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD3THSP_SD_F_SO_R 0.1
`define FD3THSP_CD_F_SO_F 0.1
`define FD3THSP_CD_R_SO_R 0.1
`define FD3THSP_CP_R_SO_R 0.1
`define FD3THSP_CP_R_SO_F 0.1
`define FD3THSP_SD_F_QN_F 0.1
`define FD3THSP_CD_F_QN_R 0.1
`define FD3THSP_CD_R_QN_F 0.1
`define FD3THSP_CP_R_QN_F 0.1
`define FD3THSP_CP_R_QN_R 0.1
`define FD3THSP_SD_F_Q_R 0.1
`define FD3THSP_CD_F_Q_F 0.1
`define FD3THSP_CD_R_Q_R 0.1
`define FD3THSP_CP_R_Q_R 0.1
`define FD3THSP_CP_R_Q_F 0.1
`define FD3THSP_CD_SD_REM_posedge_posedge 0.1
`define FD3THSP_CD_SD_REC_posedge_posedge 0.1
`define FD3THSP_CD_CP_REM_posedge_posedge 0.1
`define FD3THSP_SD_CP_REM_posedge_posedge 0.1
`define FD3THSP_CD_CP_REC_posedge_posedge 0.1
`define FD3THSP_SD_CP_REC_posedge_posedge 0.1
`define FD3THSP_CD_PWL 0.1
`define FD3THSP_SD_PWL 0.1
`define FD3THSP_CP_PWH 0.1
`define FD3THSP_CP_PWL 0.1
`define FD3THSP_D_CP_SETUP_posedge_posedge 0.1
`define FD3THSP_D_CP_SETUP_negedge_posedge 0.1
`define FD3THSP_D_CP_HOLD_posedge_posedge 0.1
`define FD3THSP_D_CP_HOLD_negedge_posedge 0.1
`define FD3THSP_TI_CP_SETUP_posedge_posedge 0.1
`define FD3THSP_TI_CP_SETUP_negedge_posedge 0.1
`define FD3THSP_TI_CP_HOLD_posedge_posedge 0.1
`define FD3THSP_TI_CP_HOLD_negedge_posedge 0.1
`define FD3THSP_TE_CP_SETUP_posedge_posedge 0.1
`define FD3THSP_TE_CP_SETUP_negedge_posedge 0.1
`define FD3THSP_TE_CP_HOLD_posedge_posedge 0.1
`define FD3THSP_TE_CP_HOLD_negedge_posedge 0.1

module FD3THSP (Q, QN, SO, D, CP, CD, SD, TI, TE);

   output Q;
   output QN;
   output SO;
   input D;
   input CP;
   input CD;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_SN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, SD, Notifier);

   buf  u2 (Q, IQ);
   buf  u3 (SO, IQ);
   not  u4 (QN, IQ);



`ifdef functional
`else
   and  (AndCDSD_, CD, SD);
   not  (TEX, TE);
   and  (AndCDSDTEX_, CD, SD, TEX);
   and  (AndCDSDTE_, CD, SD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_CDSD_, XorDTI_, CD, SD);
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);
 
   not  (D_orTI_onTE, DorTIonTE);
 
   and  (AndSDDorTI, SD, DorTIonTE);
   and  (AndCDD_orTI_, CD, D_orTI_onTE);

   specify
`ifdef verifault

      if(!TE && CD && SD) (posedge CP => (Q +: D)) = (`FD3THSP_CP_R_Q_R, `FD3THSP_CP_R_Q_F);
      if(TE && CD && SD) (posedge CP => (Q +: TI)) = (`FD3THSP_CP_R_Q_R, `FD3THSP_CP_R_Q_F);
      if(!D && TI && CD && SD) (posedge CP => (Q +: TE)) = (`FD3THSP_CP_R_Q_R, `FD3THSP_CP_R_Q_F);
      if(!TI && D && CD && SD) (posedge CP => (Q -: TE)) = (`FD3THSP_CP_R_Q_R, `FD3THSP_CP_R_Q_F);
      if(!TE && CD && SD) (posedge CP => (QN -: D)) = (`FD3THSP_CP_R_QN_R, `FD3THSP_CP_R_QN_F);
      if(TE && CD && SD) (posedge CP => (QN -: TI)) = (`FD3THSP_CP_R_QN_R, `FD3THSP_CP_R_QN_F);
      if(!D && TI && CD && SD) (posedge CP => (QN -: TE)) = (`FD3THSP_CP_R_QN_R, `FD3THSP_CP_R_QN_F);
      if(!TI && D && CD && SD) (posedge CP => (QN +: TE)) = (`FD3THSP_CP_R_QN_R, `FD3THSP_CP_R_QN_F);
      if(!TE && CD && SD) (posedge CP => (SO +: D)) = (`FD3THSP_CP_R_SO_R, `FD3THSP_CP_R_SO_F);
      if(TE && CD && SD) (posedge CP => (SO +: TI)) = (`FD3THSP_CP_R_SO_R, `FD3THSP_CP_R_SO_F);
      if(!D && TI && CD && SD) (posedge CP => (SO +: TE)) = (`FD3THSP_CP_R_SO_R, `FD3THSP_CP_R_SO_F);
      if(!TI && D && CD && SD) (posedge CP => (SO -: TE)) = (`FD3THSP_CP_R_SO_R, `FD3THSP_CP_R_SO_F);
      if(!SD) (posedge CD => (Q +: 1'b1)) = (`FD3THSP_CD_R_Q_R,`FD3THSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3THSP_CD_R_Q_R,`FD3THSP_CD_F_Q_F);
      if(CD) (negedge SD => (Q +: 1'b1)) = (`FD3THSP_SD_F_Q_R,`FD3THSP_SD_F_Q_R);
      if(!SD) (posedge CD => (QN +: 1'b0)) = (`FD3THSP_CD_F_QN_R,`FD3THSP_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`FD3THSP_CD_F_QN_R,`FD3THSP_CD_R_QN_F);
      if(CD) (negedge SD => (QN +: 1'b0)) = (`FD3THSP_SD_F_QN_F,`FD3THSP_SD_F_QN_F);
      if(!SD) (posedge CD => (SO +: 1'b1)) = (`FD3THSP_CD_R_SO_R,`FD3THSP_CD_F_SO_F);
      (negedge CD => (SO +: 1'b0)) = (`FD3THSP_CD_R_SO_R,`FD3THSP_CD_F_SO_F);
      if(CD) (negedge SD => (SO +: 1'b1)) = (`FD3THSP_SD_F_SO_R,`FD3THSP_SD_F_SO_R);

	$setuphold(posedge CP &&& AndXorDTI_CDSD_, posedge TE, `FD3THSP_TE_CP_SETUP_posedge_posedge, `FD3THSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CDSD_, negedge TE, `FD3THSP_TE_CP_SETUP_negedge_posedge, `FD3THSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDSDTE_, posedge TI, `FD3THSP_TI_CP_SETUP_posedge_posedge, `FD3THSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSDTE_, negedge TI, `FD3THSP_TI_CP_SETUP_negedge_posedge, `FD3THSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDSDTEX_, posedge D, `FD3THSP_D_CP_SETUP_posedge_posedge, `FD3THSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSDTEX_, negedge D, `FD3THSP_D_CP_SETUP_negedge_posedge, `FD3THSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD3THSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3THSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3THSP_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3THSP_CD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& AndCDD_orTI_, `FD3THSP_SD_CP_REC_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge CP &&& AndSDDorTI, `FD3THSP_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndCDD_orTI_, posedge SD, `FD3THSP_SD_CP_REM_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndSDDorTI, posedge CD, `FD3THSP_CD_CP_REM_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge SD, `FD3THSP_CD_SD_REC_posedge_posedge, Notifier);

	$hold(posedge SD, posedge CD, `FD3THSP_CD_SD_REM_posedge_posedge, Notifier);
`else

      (posedge CP => (Q +: Mux21DTITE_)) = (`FD3THSP_CP_R_Q_R, `FD3THSP_CP_R_Q_F);
      (posedge CP => (QN -: Mux21DTITE_)) = (`FD3THSP_CP_R_QN_R, `FD3THSP_CP_R_QN_F);
      (posedge CP => (SO +: Mux21DTITE_)) = (`FD3THSP_CP_R_SO_R, `FD3THSP_CP_R_SO_F);
      (posedge CD => (Q +: 1'b1)) = (`FD3THSP_CD_R_Q_R,`FD3THSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3THSP_CD_R_Q_R,`FD3THSP_CD_F_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD3THSP_SD_F_Q_R,`FD3THSP_SD_F_Q_R);
      (posedge CD => (QN +: 1'b0)) = (`FD3THSP_CD_F_QN_R,`FD3THSP_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`FD3THSP_CD_F_QN_R,`FD3THSP_CD_R_QN_F);
      (negedge SD => (QN +: 1'b0)) = (`FD3THSP_SD_F_QN_F,`FD3THSP_SD_F_QN_F);
      (posedge CD => (SO +: 1'b1)) = (`FD3THSP_CD_R_SO_R,`FD3THSP_CD_F_SO_F);
      (negedge CD => (SO +: 1'b0)) = (`FD3THSP_CD_R_SO_R,`FD3THSP_CD_F_SO_F);
      (negedge SD => (SO +: 1'b1)) = (`FD3THSP_SD_F_SO_R,`FD3THSP_SD_F_SO_R);
 
        $setuphold(posedge CP &&& AndXorDTI_CDSD_, posedge TE, `FD3THSP_TE_CP_SETUP_posedge_posedge, `FD3THSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CDSD_, negedge TE, `FD3THSP_TE_CP_SETUP_negedge_posedge, `FD3THSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDSDTE_, posedge TI, `FD3THSP_TI_CP_SETUP_posedge_posedge, `FD3THSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSDTE_, negedge TI, `FD3THSP_TI_CP_SETUP_negedge_posedge, `FD3THSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDSDTEX_, posedge D, `FD3THSP_D_CP_SETUP_posedge_posedge, `FD3THSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSDTEX_, negedge D, `FD3THSP_D_CP_SETUP_negedge_posedge, `FD3THSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD3THSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3THSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3THSP_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3THSP_CD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& AndCDD_orTI_, `FD3THSP_SD_CP_REC_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge CP &&& AndSDDorTI, `FD3THSP_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndCDD_orTI_, posedge SD, `FD3THSP_SD_CP_REM_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndSDDorTI, posedge CD, `FD3THSP_CD_CP_REM_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge SD, `FD3THSP_CD_SD_REC_posedge_posedge, Notifier);
 
        $hold(posedge SD, posedge CD, `FD3THSP_CD_SD_REM_posedge_posedge, Notifier);
`endif

   endspecify
`endif


endmodule // FD3THSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:11 and Version :1.1 //
 
//  START 
// CELL FD3TQHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD3TQHS_SD_F_SO_R 0.1
`define FD3TQHS_CD_F_SO_F 0.1
`define FD3TQHS_CD_R_SO_R 0.1
`define FD3TQHS_CP_R_SO_R 0.1
`define FD3TQHS_CP_R_SO_F 0.1
`define FD3TQHS_SD_F_Q_R 0.1
`define FD3TQHS_CD_F_Q_F 0.1
`define FD3TQHS_CD_R_Q_R 0.1
`define FD3TQHS_CP_R_Q_R 0.1
`define FD3TQHS_CP_R_Q_F 0.1
`define FD3TQHS_CD_SD_REM_posedge_posedge 0.1
`define FD3TQHS_CD_SD_REC_posedge_posedge 0.1
`define FD3TQHS_CD_CP_REM_posedge_posedge 0.1
`define FD3TQHS_SD_CP_REM_posedge_posedge 0.1
`define FD3TQHS_CD_CP_REC_posedge_posedge 0.1
`define FD3TQHS_SD_CP_REC_posedge_posedge 0.1
`define FD3TQHS_CD_PWL 0.1
`define FD3TQHS_SD_PWL 0.1
`define FD3TQHS_CP_PWH 0.1
`define FD3TQHS_CP_PWL 0.1
`define FD3TQHS_D_CP_SETUP_posedge_posedge 0.1
`define FD3TQHS_D_CP_SETUP_negedge_posedge 0.1
`define FD3TQHS_D_CP_HOLD_posedge_posedge 0.1
`define FD3TQHS_D_CP_HOLD_negedge_posedge 0.1
`define FD3TQHS_TI_CP_SETUP_posedge_posedge 0.1
`define FD3TQHS_TI_CP_SETUP_negedge_posedge 0.1
`define FD3TQHS_TI_CP_HOLD_posedge_posedge 0.1
`define FD3TQHS_TI_CP_HOLD_negedge_posedge 0.1
`define FD3TQHS_TE_CP_SETUP_posedge_posedge 0.1
`define FD3TQHS_TE_CP_SETUP_negedge_posedge 0.1
`define FD3TQHS_TE_CP_HOLD_posedge_posedge 0.1
`define FD3TQHS_TE_CP_HOLD_negedge_posedge 0.1

module FD3TQHS (Q, SO, D, CP, CD, SD, TI, TE);

   output Q;
   output SO;
   input D;
   input CP;
   input CD;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_SN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, SD, Notifier);

   buf  u2 (Q, IQ);
   buf  u3 (SO, IQ);



`ifdef functional
`else
   and  (AndCDSD_, CD, SD);
   not  (TEX, TE);
   and  (AndCDSDTEX_, CD, SD, TEX);
   and  (AndCDSDTE_, CD, SD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_CDSD_, XorDTI_, CD, SD);
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);
 
   not  (D_orTI_onTE, DorTIonTE);
 
   and  (AndSDDorTI, SD, DorTIonTE);
   and  (AndCDD_orTI_, CD, D_orTI_onTE);

   specify
`ifdef verifault
      if(!TE && CD && SD) (posedge CP => (Q +: D)) = (`FD3TQHS_CP_R_Q_R, `FD3TQHS_CP_R_Q_F);
      if(TE && CD && SD) (posedge CP => (Q +: TI)) = (`FD3TQHS_CP_R_Q_R, `FD3TQHS_CP_R_Q_F);
      if(!D && TI && CD && SD) (posedge CP => (Q +: TE)) = (`FD3TQHS_CP_R_Q_R, `FD3TQHS_CP_R_Q_F);
      if(!TI && D && CD && SD) (posedge CP => (Q -: TE)) = (`FD3TQHS_CP_R_Q_R, `FD3TQHS_CP_R_Q_F);
      if(!TE && CD && SD) (posedge CP => (SO +: D)) = (`FD3TQHS_CP_R_SO_R, `FD3TQHS_CP_R_SO_F);
      if(TE && CD && SD) (posedge CP => (SO +: TI)) = (`FD3TQHS_CP_R_SO_R, `FD3TQHS_CP_R_SO_F);
      if(!D && TI && CD && SD) (posedge CP => (SO +: TE)) = (`FD3TQHS_CP_R_SO_R, `FD3TQHS_CP_R_SO_F);
      if(!TI && D && CD && SD) (posedge CP => (SO -: TE)) = (`FD3TQHS_CP_R_SO_R, `FD3TQHS_CP_R_SO_F);
      if(!SD) (posedge CD => (Q +: 1'b1)) = (`FD3TQHS_CD_R_Q_R,`FD3TQHS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3TQHS_CD_R_Q_R,`FD3TQHS_CD_F_Q_F);
      if(CD) (negedge SD => (Q +: 1'b1)) = (`FD3TQHS_SD_F_Q_R,`FD3TQHS_SD_F_Q_R);
      if(!SD) (posedge CD => (SO +: 1'b1)) = (`FD3TQHS_CD_R_SO_R,`FD3TQHS_CD_F_SO_F);
      (negedge CD => (SO +: 1'b0)) = (`FD3TQHS_CD_R_SO_R,`FD3TQHS_CD_F_SO_F);
      if(CD) (negedge SD => (SO +: 1'b1)) = (`FD3TQHS_SD_F_SO_R,`FD3TQHS_SD_F_SO_R);

	$setuphold(posedge CP &&& AndXorDTI_CDSD_, posedge TE, `FD3TQHS_TE_CP_SETUP_posedge_posedge, `FD3TQHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CDSD_, negedge TE, `FD3TQHS_TE_CP_SETUP_negedge_posedge, `FD3TQHS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDSDTE_, posedge TI, `FD3TQHS_TI_CP_SETUP_posedge_posedge, `FD3TQHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSDTE_, negedge TI, `FD3TQHS_TI_CP_SETUP_negedge_posedge, `FD3TQHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDSDTEX_, posedge D, `FD3TQHS_D_CP_SETUP_posedge_posedge, `FD3TQHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSDTEX_, negedge D, `FD3TQHS_D_CP_SETUP_negedge_posedge, `FD3TQHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD3TQHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3TQHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3TQHS_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3TQHS_CD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& AndCDD_orTI_, `FD3TQHS_SD_CP_REC_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge CP &&& AndSDDorTI, `FD3TQHS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndCDD_orTI_, posedge SD, `FD3TQHS_SD_CP_REM_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndSDDorTI, posedge CD, `FD3TQHS_CD_CP_REM_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge SD, `FD3TQHS_CD_SD_REC_posedge_posedge, Notifier);

	$hold(posedge SD, posedge CD, `FD3TQHS_CD_SD_REM_posedge_posedge, Notifier);

`else 
      (posedge CP => (Q +: Mux21DTITE_)) = (`FD3TQHS_CP_R_Q_R, `FD3TQHS_CP_R_Q_F);
      (posedge CP => (SO +: Mux21DTITE_)) = (`FD3TQHS_CP_R_SO_R, `FD3TQHS_CP_R_SO_F);
      (posedge CD => (Q +: 1'b1)) = (`FD3TQHS_CD_R_Q_R,`FD3TQHS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3TQHS_CD_R_Q_R,`FD3TQHS_CD_F_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD3TQHS_SD_F_Q_R,`FD3TQHS_SD_F_Q_R);
      (posedge CD => (SO +: 1'b1)) = (`FD3TQHS_CD_R_SO_R,`FD3TQHS_CD_F_SO_F);
      (negedge CD => (SO +: 1'b0)) = (`FD3TQHS_CD_R_SO_R,`FD3TQHS_CD_F_SO_F);
      (negedge SD => (SO +: 1'b1)) = (`FD3TQHS_SD_F_SO_R,`FD3TQHS_SD_F_SO_R);
 
        $setuphold(posedge CP &&& AndXorDTI_CDSD_, posedge TE, `FD3TQHS_TE_CP_SETUP_posedge_posedge, `FD3TQHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CDSD_, negedge TE, `FD3TQHS_TE_CP_SETUP_negedge_posedge, `FD3TQHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDSDTE_, posedge TI, `FD3TQHS_TI_CP_SETUP_posedge_posedge, `FD3TQHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSDTE_, negedge TI, `FD3TQHS_TI_CP_SETUP_negedge_posedge, `FD3TQHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDSDTEX_, posedge D, `FD3TQHS_D_CP_SETUP_posedge_posedge, `FD3TQHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSDTEX_, negedge D, `FD3TQHS_D_CP_SETUP_negedge_posedge, `FD3TQHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD3TQHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3TQHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3TQHS_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3TQHS_CD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& AndCDD_orTI_, `FD3TQHS_SD_CP_REC_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge CP &&& AndSDDorTI, `FD3TQHS_CD_CP_REC_posedge_posedge,Notifier);
        $hold(posedge CP &&& AndCDD_orTI_, posedge SD, `FD3TQHS_SD_CP_REM_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndSDDorTI, posedge CD, `FD3TQHS_CD_CP_REM_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge SD, `FD3TQHS_CD_SD_REC_posedge_posedge, Notifier);
 
        $hold(posedge SD, posedge CD, `FD3TQHS_CD_SD_REM_posedge_posedge, Notifier);
 
`endif 

   endspecify
`endif


endmodule // FD3TQHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:15 and Version :1.1 //
 
//  START 
// CELL FD3TQHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD3TQHSP_SD_F_SO_R 0.1
`define FD3TQHSP_CD_F_SO_F 0.1
`define FD3TQHSP_CD_R_SO_R 0.1
`define FD3TQHSP_CP_R_SO_R 0.1
`define FD3TQHSP_CP_R_SO_F 0.1
`define FD3TQHSP_SD_F_Q_R 0.1
`define FD3TQHSP_CD_F_Q_F 0.1
`define FD3TQHSP_CD_R_Q_R 0.1
`define FD3TQHSP_CP_R_Q_R 0.1
`define FD3TQHSP_CP_R_Q_F 0.1
`define FD3TQHSP_CD_SD_REM_posedge_posedge 0.1
`define FD3TQHSP_CD_SD_REC_posedge_posedge 0.1
`define FD3TQHSP_CD_CP_REM_posedge_posedge 0.1
`define FD3TQHSP_SD_CP_REM_posedge_posedge 0.1
`define FD3TQHSP_CD_CP_REC_posedge_posedge 0.1
`define FD3TQHSP_SD_CP_REC_posedge_posedge 0.1
`define FD3TQHSP_CD_PWL 0.1
`define FD3TQHSP_SD_PWL 0.1
`define FD3TQHSP_CP_PWH 0.1
`define FD3TQHSP_CP_PWL 0.1
`define FD3TQHSP_D_CP_SETUP_posedge_posedge 0.1
`define FD3TQHSP_D_CP_SETUP_negedge_posedge 0.1
`define FD3TQHSP_D_CP_HOLD_posedge_posedge 0.1
`define FD3TQHSP_D_CP_HOLD_negedge_posedge 0.1
`define FD3TQHSP_TI_CP_SETUP_posedge_posedge 0.1
`define FD3TQHSP_TI_CP_SETUP_negedge_posedge 0.1
`define FD3TQHSP_TI_CP_HOLD_posedge_posedge 0.1
`define FD3TQHSP_TI_CP_HOLD_negedge_posedge 0.1
`define FD3TQHSP_TE_CP_SETUP_posedge_posedge 0.1
`define FD3TQHSP_TE_CP_SETUP_negedge_posedge 0.1
`define FD3TQHSP_TE_CP_HOLD_posedge_posedge 0.1
`define FD3TQHSP_TE_CP_HOLD_negedge_posedge 0.1

module FD3TQHSP (Q, SO, D, CP, CD, SD, TI, TE);

   output Q;
   output SO;
   input D;
   input CP;
   input CD;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_SN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, SD, Notifier);

   buf  u2 (Q, IQ);
   buf  u3 (SO, IQ);



`ifdef functional
`else
   and  (AndCDSD_, CD, SD);
   not  (TEX, TE);
   and  (AndCDSDTEX_, CD, SD, TEX);
   and  (AndCDSDTE_, CD, SD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_CDSD_, XorDTI_, CD, SD);
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);
 
   not  (D_orTI_onTE, DorTIonTE);
 
   and  (AndSDDorTI, SD, DorTIonTE);
   and  (AndCDD_orTI_, CD, D_orTI_onTE);

   specify
`ifdef verifault
      if(!TE && CD && SD) (posedge CP => (Q +: D)) = (`FD3TQHSP_CP_R_Q_R, `FD3TQHSP_CP_R_Q_F);
      if(TE && CD && SD) (posedge CP => (Q +: TI)) = (`FD3TQHSP_CP_R_Q_R, `FD3TQHSP_CP_R_Q_F);
      if(!D && TI && CD && SD) (posedge CP => (Q +: TE)) = (`FD3TQHSP_CP_R_Q_R, `FD3TQHSP_CP_R_Q_F);
      if(!TI && D && CD && SD) (posedge CP => (Q -: TE)) = (`FD3TQHSP_CP_R_Q_R, `FD3TQHSP_CP_R_Q_F);
      if(!TE && CD && SD) (posedge CP => (SO +: D)) = (`FD3TQHSP_CP_R_SO_R, `FD3TQHSP_CP_R_SO_F);
      if(TE && CD && SD) (posedge CP => (SO +: TI)) = (`FD3TQHSP_CP_R_SO_R, `FD3TQHSP_CP_R_SO_F);
      if(!D && TI && CD && SD) (posedge CP => (SO +: TE)) = (`FD3TQHSP_CP_R_SO_R, `FD3TQHSP_CP_R_SO_F);
      if(!TI && D && CD && SD) (posedge CP => (SO -: TE)) = (`FD3TQHSP_CP_R_SO_R, `FD3TQHSP_CP_R_SO_F);
      if(!SD) (posedge CD => (Q +: 1'b1)) = (`FD3TQHSP_CD_R_Q_R,`FD3TQHSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3TQHSP_CD_R_Q_R,`FD3TQHSP_CD_F_Q_F);
      if(CD) (negedge SD => (Q +: 1'b1)) = (`FD3TQHSP_SD_F_Q_R,`FD3TQHSP_SD_F_Q_R);
      if(!SD) (posedge CD => (SO +: 1'b1)) = (`FD3TQHSP_CD_R_SO_R,`FD3TQHSP_CD_F_SO_F);
      (negedge CD => (SO +: 1'b0)) = (`FD3TQHSP_CD_R_SO_R,`FD3TQHSP_CD_F_SO_F);
      if(CD) (negedge SD => (SO +: 1'b1)) = (`FD3TQHSP_SD_F_SO_R,`FD3TQHSP_SD_F_SO_R);

	$setuphold(posedge CP &&& AndXorDTI_CDSD_, posedge TE, `FD3TQHSP_TE_CP_SETUP_posedge_posedge, `FD3TQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CDSD_, negedge TE, `FD3TQHSP_TE_CP_SETUP_negedge_posedge, `FD3TQHSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDSDTE_, posedge TI, `FD3TQHSP_TI_CP_SETUP_posedge_posedge, `FD3TQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSDTE_, negedge TI, `FD3TQHSP_TI_CP_SETUP_negedge_posedge, `FD3TQHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDSDTEX_, posedge D, `FD3TQHSP_D_CP_SETUP_posedge_posedge, `FD3TQHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSDTEX_, negedge D, `FD3TQHSP_D_CP_SETUP_negedge_posedge, `FD3TQHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD3TQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3TQHSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3TQHSP_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3TQHSP_CD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& AndCDD_orTI_, `FD3TQHSP_SD_CP_REC_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge CP &&& AndSDDorTI, `FD3TQHSP_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndCDD_orTI_, posedge SD, `FD3TQHSP_SD_CP_REM_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndSDDorTI, posedge CD, `FD3TQHSP_CD_CP_REM_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge SD, `FD3TQHSP_CD_SD_REC_posedge_posedge, Notifier);

	$hold(posedge SD, posedge CD, `FD3TQHSP_CD_SD_REM_posedge_posedge, Notifier);

`else 
      (posedge CP => (Q +: Mux21DTITE_)) = (`FD3TQHSP_CP_R_Q_R, `FD3TQHSP_CP_R_Q_F);
      (posedge CP => (SO +: Mux21DTITE_)) = (`FD3TQHSP_CP_R_SO_R, `FD3TQHSP_CP_R_SO_F);
      (posedge CD => (Q +: 1'b1)) = (`FD3TQHSP_CD_R_Q_R,`FD3TQHSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3TQHSP_CD_R_Q_R,`FD3TQHSP_CD_F_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD3TQHSP_SD_F_Q_R,`FD3TQHSP_SD_F_Q_R);
      (posedge CD => (SO +: 1'b1)) = (`FD3TQHSP_CD_R_SO_R,`FD3TQHSP_CD_F_SO_F);
      (negedge CD => (SO +: 1'b0)) = (`FD3TQHSP_CD_R_SO_R,`FD3TQHSP_CD_F_SO_F);
      (negedge SD => (SO +: 1'b1)) = (`FD3TQHSP_SD_F_SO_R,`FD3TQHSP_SD_F_SO_R);
 
        $setuphold(posedge CP &&& AndXorDTI_CDSD_, posedge TE, `FD3TQHSP_TE_CP_SETUP_posedge_posedge, `FD3TQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CDSD_, negedge TE, `FD3TQHSP_TE_CP_SETUP_negedge_posedge, `FD3TQHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDSDTE_, posedge TI, `FD3TQHSP_TI_CP_SETUP_posedge_posedge, `FD3TQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSDTE_, negedge TI, `FD3TQHSP_TI_CP_SETUP_negedge_posedge, `FD3TQHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDSDTEX_, posedge D, `FD3TQHSP_D_CP_SETUP_posedge_posedge, `FD3TQHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSDTEX_, negedge D, `FD3TQHSP_D_CP_SETUP_negedge_posedge, `FD3TQHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD3TQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3TQHSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3TQHSP_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3TQHSP_CD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& AndCDD_orTI_, `FD3TQHSP_SD_CP_REC_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge CP &&& AndSDDorTI, `FD3TQHSP_CD_CP_REC_posedge_posedge,Notifier);
        $hold(posedge CP &&& AndCDD_orTI_, posedge SD, `FD3TQHSP_SD_CP_REM_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndSDDorTI, posedge CD, `FD3TQHSP_CD_CP_REM_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge SD, `FD3TQHSP_CD_SD_REC_posedge_posedge, Notifier);
 
        $hold(posedge SD, posedge CD, `FD3TQHSP_CD_SD_REM_posedge_posedge, Notifier);
 
`endif 

   endspecify
`endif


endmodule // FD3TQHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:15 and Version :1.1 //
 
//  START 
// CELL FD3TQHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD3TQHSX4_SD_F_SO_R 0.1
`define FD3TQHSX4_CD_F_SO_F 0.1
`define FD3TQHSX4_CD_R_SO_R 0.1
`define FD3TQHSX4_CP_R_SO_R 0.1
`define FD3TQHSX4_CP_R_SO_F 0.1
`define FD3TQHSX4_SD_F_Q_R 0.1
`define FD3TQHSX4_CD_F_Q_F 0.1
`define FD3TQHSX4_CD_R_Q_R 0.1
`define FD3TQHSX4_CP_R_Q_R 0.1
`define FD3TQHSX4_CP_R_Q_F 0.1
`define FD3TQHSX4_CD_SD_REM_posedge_posedge 0.1
`define FD3TQHSX4_CD_SD_REC_posedge_posedge 0.1
`define FD3TQHSX4_CD_CP_REM_posedge_posedge 0.1
`define FD3TQHSX4_SD_CP_REM_posedge_posedge 0.1
`define FD3TQHSX4_CD_CP_REC_posedge_posedge 0.1
`define FD3TQHSX4_SD_CP_REC_posedge_posedge 0.1
`define FD3TQHSX4_CD_PWL 0.1
`define FD3TQHSX4_SD_PWL 0.1
`define FD3TQHSX4_CP_PWH 0.1
`define FD3TQHSX4_CP_PWL 0.1
`define FD3TQHSX4_D_CP_SETUP_posedge_posedge 0.1
`define FD3TQHSX4_D_CP_SETUP_negedge_posedge 0.1
`define FD3TQHSX4_D_CP_HOLD_posedge_posedge 0.1
`define FD3TQHSX4_D_CP_HOLD_negedge_posedge 0.1
`define FD3TQHSX4_TI_CP_SETUP_posedge_posedge 0.1
`define FD3TQHSX4_TI_CP_SETUP_negedge_posedge 0.1
`define FD3TQHSX4_TI_CP_HOLD_posedge_posedge 0.1
`define FD3TQHSX4_TI_CP_HOLD_negedge_posedge 0.1
`define FD3TQHSX4_TE_CP_SETUP_posedge_posedge 0.1
`define FD3TQHSX4_TE_CP_SETUP_negedge_posedge 0.1
`define FD3TQHSX4_TE_CP_HOLD_posedge_posedge 0.1
`define FD3TQHSX4_TE_CP_HOLD_negedge_posedge 0.1

module FD3TQHSX4 (Q, SO, D, CP, CD, SD, TI, TE);

   output Q;
   output SO;
   input D;
   input CP;
   input CD;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_RN_SN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, CD, SD, Notifier);

   buf  u2 (Q, IQ);
   buf  u3 (SO, IQ);



`ifdef functional
`else
   and  (AndCDSD_, CD, SD);
   not  (TEX, TE);
   and  (AndCDSDTEX_, CD, SD, TEX);
   and  (AndCDSDTE_, CD, SD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_CDSD_, XorDTI_, CD, SD);
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);
 
   not  (D_orTI_onTE, DorTIonTE);
 
   and  (AndSDDorTI, SD, DorTIonTE);
   and  (AndCDD_orTI_, CD, D_orTI_onTE);

   specify
`ifdef verifault
      if(!TE && CD && SD) (posedge CP => (Q +: D)) = (`FD3TQHSX4_CP_R_Q_R, `FD3TQHSX4_CP_R_Q_F);
      if(TE && CD && SD) (posedge CP => (Q +: TI)) = (`FD3TQHSX4_CP_R_Q_R, `FD3TQHSX4_CP_R_Q_F);
      if(!D && TI && CD && SD) (posedge CP => (Q +: TE)) = (`FD3TQHSX4_CP_R_Q_R, `FD3TQHSX4_CP_R_Q_F);
      if(!TI && D && CD && SD) (posedge CP => (Q -: TE)) = (`FD3TQHSX4_CP_R_Q_R, `FD3TQHSX4_CP_R_Q_F);
      if(!TE && CD && SD) (posedge CP => (SO +: D)) = (`FD3TQHSX4_CP_R_SO_R, `FD3TQHSX4_CP_R_SO_F);
      if(TE && CD && SD) (posedge CP => (SO +: TI)) = (`FD3TQHSX4_CP_R_SO_R, `FD3TQHSX4_CP_R_SO_F);
      if(!D && TI && CD && SD) (posedge CP => (SO +: TE)) = (`FD3TQHSX4_CP_R_SO_R, `FD3TQHSX4_CP_R_SO_F);
      if(!TI && D && CD && SD) (posedge CP => (SO -: TE)) = (`FD3TQHSX4_CP_R_SO_R, `FD3TQHSX4_CP_R_SO_F);
      if(!SD) (posedge CD => (Q +: 1'b1)) = (`FD3TQHSX4_CD_R_Q_R,`FD3TQHSX4_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3TQHSX4_CD_R_Q_R,`FD3TQHSX4_CD_F_Q_F);
      if(CD) (negedge SD => (Q +: 1'b1)) = (`FD3TQHSX4_SD_F_Q_R,`FD3TQHSX4_SD_F_Q_R);
      if(!SD) (posedge CD => (SO +: 1'b1)) = (`FD3TQHSX4_CD_R_SO_R,`FD3TQHSX4_CD_F_SO_F);
      (negedge CD => (SO +: 1'b0)) = (`FD3TQHSX4_CD_R_SO_R,`FD3TQHSX4_CD_F_SO_F);
      if(CD) (negedge SD => (SO +: 1'b1)) = (`FD3TQHSX4_SD_F_SO_R,`FD3TQHSX4_SD_F_SO_R);

	$setuphold(posedge CP &&& AndXorDTI_CDSD_, posedge TE, `FD3TQHSX4_TE_CP_SETUP_posedge_posedge, `FD3TQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_CDSD_, negedge TE, `FD3TQHSX4_TE_CP_SETUP_negedge_posedge, `FD3TQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDSDTE_, posedge TI, `FD3TQHSX4_TI_CP_SETUP_posedge_posedge, `FD3TQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSDTE_, negedge TI, `FD3TQHSX4_TI_CP_SETUP_negedge_posedge, `FD3TQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDSDTEX_, posedge D, `FD3TQHSX4_D_CP_SETUP_posedge_posedge, `FD3TQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSDTEX_, negedge D, `FD3TQHSX4_D_CP_SETUP_negedge_posedge, `FD3TQHSX4_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD3TQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3TQHSX4_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3TQHSX4_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3TQHSX4_CD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& AndCDD_orTI_, `FD3TQHSX4_SD_CP_REC_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge CP &&& AndSDDorTI, `FD3TQHSX4_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndCDD_orTI_, posedge SD, `FD3TQHSX4_SD_CP_REM_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndSDDorTI, posedge CD, `FD3TQHSX4_CD_CP_REM_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge SD, `FD3TQHSX4_CD_SD_REC_posedge_posedge, Notifier);

	$hold(posedge SD, posedge CD, `FD3TQHSX4_CD_SD_REM_posedge_posedge, Notifier);

`else 
      (posedge CP => (Q +: Mux21DTITE_)) = (`FD3TQHSX4_CP_R_Q_R, `FD3TQHSX4_CP_R_Q_F);
      (posedge CP => (SO +: Mux21DTITE_)) = (`FD3TQHSX4_CP_R_SO_R, `FD3TQHSX4_CP_R_SO_F);
      (posedge CD => (Q +: 1'b1)) = (`FD3TQHSX4_CD_R_Q_R,`FD3TQHSX4_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FD3TQHSX4_CD_R_Q_R,`FD3TQHSX4_CD_F_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD3TQHSX4_SD_F_Q_R,`FD3TQHSX4_SD_F_Q_R);
      (posedge CD => (SO +: 1'b1)) = (`FD3TQHSX4_CD_R_SO_R,`FD3TQHSX4_CD_F_SO_F);
      (negedge CD => (SO +: 1'b0)) = (`FD3TQHSX4_CD_R_SO_R,`FD3TQHSX4_CD_F_SO_F);
      (negedge SD => (SO +: 1'b1)) = (`FD3TQHSX4_SD_F_SO_R,`FD3TQHSX4_SD_F_SO_R);
 
        $setuphold(posedge CP &&& AndXorDTI_CDSD_, posedge TE, `FD3TQHSX4_TE_CP_SETUP_posedge_posedge, `FD3TQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_CDSD_, negedge TE, `FD3TQHSX4_TE_CP_SETUP_negedge_posedge, `FD3TQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDSDTE_, posedge TI, `FD3TQHSX4_TI_CP_SETUP_posedge_posedge, `FD3TQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSDTE_, negedge TI, `FD3TQHSX4_TI_CP_SETUP_negedge_posedge, `FD3TQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDSDTEX_, posedge D, `FD3TQHSX4_D_CP_SETUP_posedge_posedge, `FD3TQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSDTEX_, negedge D, `FD3TQHSX4_D_CP_SETUP_negedge_posedge, `FD3TQHSX4_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD3TQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FD3TQHSX4_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD3TQHSX4_SD_PWL, 0, Notifier);
      $width(negedge CD, `FD3TQHSX4_CD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& AndCDD_orTI_, `FD3TQHSX4_SD_CP_REC_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge CP &&& AndSDDorTI, `FD3TQHSX4_CD_CP_REC_posedge_posedge,Notifier);
        $hold(posedge CP &&& AndCDD_orTI_, posedge SD, `FD3TQHSX4_SD_CP_REM_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndSDDorTI, posedge CD, `FD3TQHSX4_CD_CP_REM_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge SD, `FD3TQHSX4_CD_SD_REC_posedge_posedge, Notifier);
 
        $hold(posedge SD, posedge CD, `FD3TQHSX4_CD_SD_REM_posedge_posedge, Notifier);
 
`endif 

   endspecify
`endif


endmodule // FD3TQHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:15 and Version :1.1 //
 
//  START 
// CELL FD4HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD4HS_SD_F_QN_F 0.1
`define FD4HS_CP_R_QN_F 0.1
`define FD4HS_CP_R_QN_R 0.1
`define FD4HS_SD_F_Q_R 0.1
`define FD4HS_CP_R_Q_R 0.1
`define FD4HS_CP_R_Q_F 0.1
`define FD4HS_SD_CP_REM_posedge_posedge 0.1
`define FD4HS_SD_CP_REC_posedge_posedge 0.1
`define FD4HS_SD_PWL 0.1
`define FD4HS_CP_PWH 0.1
`define FD4HS_CP_PWL 0.1
`define FD4HS_D_CP_SETUP_posedge_posedge 0.1
`define FD4HS_D_CP_SETUP_negedge_posedge 0.1
`define FD4HS_D_CP_HOLD_posedge_posedge 0.1
`define FD4HS_D_CP_HOLD_negedge_posedge 0.1

module FD4HS (Q, QN, D, CP, SD);

   output Q;
   output QN;
   input D;
   input CP;
   input SD;


   reg Notifier;


   U_FD_P_SN_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, SD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   not  (D_, D);

   specify
`ifdef verifault

      if(SD) (posedge CP => (Q +: D)) = (`FD4HS_CP_R_Q_R, `FD4HS_CP_R_Q_F);
      if(SD) (posedge CP => (QN -: D)) = (`FD4HS_CP_R_QN_R, `FD4HS_CP_R_QN_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4HS_SD_F_Q_R,`FD4HS_SD_F_Q_R);
      (negedge SD => (QN +: 1'b0)) = (`FD4HS_SD_F_QN_F,`FD4HS_SD_F_QN_F);

	$setuphold(posedge CP &&& SD, posedge D, `FD4HS_D_CP_SETUP_posedge_posedge, `FD4HS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& SD, negedge D, `FD4HS_D_CP_SETUP_negedge_posedge, `FD4HS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD4HS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4HS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4HS_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_, `FD4HS_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_, posedge SD, `FD4HS_SD_CP_REM_posedge_posedge, Notifier);


`else
      (posedge CP => (Q +: D)) = (`FD4HS_CP_R_Q_R, `FD4HS_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`FD4HS_CP_R_QN_R, `FD4HS_CP_R_QN_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4HS_SD_F_Q_R,`FD4HS_SD_F_Q_R);
      (negedge SD => (QN +: 1'b0)) = (`FD4HS_SD_F_QN_F,`FD4HS_SD_F_QN_F);
 
        $setuphold(posedge CP &&& SD, posedge D, `FD4HS_D_CP_SETUP_posedge_posedge, `FD4HS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& SD, negedge D, `FD4HS_D_CP_SETUP_negedge_posedge, `FD4HS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD4HS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4HS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4HS_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_, `FD4HS_SD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D_, posedge SD, `FD4HS_SD_CP_REM_posedge_posedge, Notifier);
 
`endif
   endspecify
`endif


endmodule // FD4HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:17 and Version :1.1 //
 
//  START 
// CELL FD4HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD4HSP_SD_F_QN_F 0.1
`define FD4HSP_CP_R_QN_F 0.1
`define FD4HSP_CP_R_QN_R 0.1
`define FD4HSP_SD_F_Q_R 0.1
`define FD4HSP_CP_R_Q_R 0.1
`define FD4HSP_CP_R_Q_F 0.1
`define FD4HSP_SD_CP_REM_posedge_posedge 0.1
`define FD4HSP_SD_CP_REC_posedge_posedge 0.1
`define FD4HSP_SD_PWL 0.1
`define FD4HSP_CP_PWH 0.1
`define FD4HSP_CP_PWL 0.1
`define FD4HSP_D_CP_SETUP_posedge_posedge 0.1
`define FD4HSP_D_CP_SETUP_negedge_posedge 0.1
`define FD4HSP_D_CP_HOLD_posedge_posedge 0.1
`define FD4HSP_D_CP_HOLD_negedge_posedge 0.1

module FD4HSP (Q, QN, D, CP, SD);

   output Q;
   output QN;
   input D;
   input CP;
   input SD;


   reg Notifier;


   U_FD_P_SN_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, SD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   not  (D_, D);

   specify
`ifdef verifault

      if(SD) (posedge CP => (Q +: D)) = (`FD4HSP_CP_R_Q_R, `FD4HSP_CP_R_Q_F);
      if(SD) (posedge CP => (QN -: D)) = (`FD4HSP_CP_R_QN_R, `FD4HSP_CP_R_QN_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4HSP_SD_F_Q_R,`FD4HSP_SD_F_Q_R);
      (negedge SD => (QN +: 1'b0)) = (`FD4HSP_SD_F_QN_F,`FD4HSP_SD_F_QN_F);

	$setuphold(posedge CP &&& SD, posedge D, `FD4HSP_D_CP_SETUP_posedge_posedge, `FD4HSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& SD, negedge D, `FD4HSP_D_CP_SETUP_negedge_posedge, `FD4HSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD4HSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4HSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4HSP_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_, `FD4HSP_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_, posedge SD, `FD4HSP_SD_CP_REM_posedge_posedge, Notifier);


`else
      (posedge CP => (Q +: D)) = (`FD4HSP_CP_R_Q_R, `FD4HSP_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`FD4HSP_CP_R_QN_R, `FD4HSP_CP_R_QN_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4HSP_SD_F_Q_R,`FD4HSP_SD_F_Q_R);
      (negedge SD => (QN +: 1'b0)) = (`FD4HSP_SD_F_QN_F,`FD4HSP_SD_F_QN_F);
 
        $setuphold(posedge CP &&& SD, posedge D, `FD4HSP_D_CP_SETUP_posedge_posedge, `FD4HSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& SD, negedge D, `FD4HSP_D_CP_SETUP_negedge_posedge, `FD4HSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD4HSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4HSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4HSP_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_, `FD4HSP_SD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D_, posedge SD, `FD4HSP_SD_CP_REM_posedge_posedge, Notifier);
 
`endif
   endspecify
`endif


endmodule // FD4HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:17 and Version :1.1 //
 
//  START 
// CELL FDM4HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDM4HS_SD_F_QN_F 0.1
`define FDM4HS_CP_R_QN_F 0.1
`define FDM4HS_CP_R_QN_R 0.1
`define FDM4HS_SD_F_Q_R 0.1
`define FDM4HS_CP_R_Q_R 0.1
`define FDM4HS_CP_R_Q_F 0.1
`define FDM4HS_SD_CP_REM_posedge_posedge 0.1
`define FDM4HS_SD_CP_REC_posedge_posedge 0.1
`define FDM4HS_SD_PWL 0.1
`define FDM4HS_CP_PWH 0.1
`define FDM4HS_CP_PWL 0.1
`define FDM4HS_D_CP_SETUP_posedge_posedge 0.1
`define FDM4HS_D_CP_SETUP_negedge_posedge 0.1
`define FDM4HS_D_CP_HOLD_posedge_posedge 0.1
`define FDM4HS_D_CP_HOLD_negedge_posedge 0.1

module FDM4HS (Q, QN, D, CP, SD);

   output Q;
   output QN;
   input D;
   input CP;
   input SD;


   reg Notifier;


   U_FD_P_SN_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, SD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   not  (D_, D);

   specify
`ifdef verifault

      if(SD) (posedge CP => (Q +: D)) = (`FDM4HS_CP_R_Q_R, `FDM4HS_CP_R_Q_F);
      if(SD) (posedge CP => (QN -: D)) = (`FDM4HS_CP_R_QN_R, `FDM4HS_CP_R_QN_F);
      (negedge SD => (Q +: 1'b1)) = (`FDM4HS_SD_F_Q_R,`FDM4HS_SD_F_Q_R);
      (negedge SD => (QN +: 1'b0)) = (`FDM4HS_SD_F_QN_F,`FDM4HS_SD_F_QN_F);

	$setuphold(posedge CP &&& SD, posedge D, `FDM4HS_D_CP_SETUP_posedge_posedge, `FDM4HS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& SD, negedge D, `FDM4HS_D_CP_SETUP_negedge_posedge, `FDM4HS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDM4HS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FDM4HS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FDM4HS_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_, `FDM4HS_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_, posedge SD, `FDM4HS_SD_CP_REM_posedge_posedge, Notifier);


`else
      (posedge CP => (Q +: D)) = (`FDM4HS_CP_R_Q_R, `FDM4HS_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`FDM4HS_CP_R_QN_R, `FDM4HS_CP_R_QN_F);
      (negedge SD => (Q +: 1'b1)) = (`FDM4HS_SD_F_Q_R,`FDM4HS_SD_F_Q_R);
      (negedge SD => (QN +: 1'b0)) = (`FDM4HS_SD_F_QN_F,`FDM4HS_SD_F_QN_F);
 
        $setuphold(posedge CP &&& SD, posedge D, `FDM4HS_D_CP_SETUP_posedge_posedge, `FDM4HS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& SD, negedge D, `FDM4HS_D_CP_SETUP_negedge_posedge, `FDM4HS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDM4HS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FDM4HS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FDM4HS_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_, `FDM4HS_SD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D_, posedge SD, `FDM4HS_SD_CP_REM_posedge_posedge, Notifier);
 
`endif
   endspecify
`endif


endmodule // FDM4HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:17 and Version :1.1 //
 
//  START 
// CELL FDM4HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDM4HSP_SD_F_QN_F 0.1
`define FDM4HSP_CP_R_QN_F 0.1
`define FDM4HSP_CP_R_QN_R 0.1
`define FDM4HSP_SD_F_Q_R 0.1
`define FDM4HSP_CP_R_Q_R 0.1
`define FDM4HSP_CP_R_Q_F 0.1
`define FDM4HSP_SD_CP_REM_posedge_posedge 0.1
`define FDM4HSP_SD_CP_REC_posedge_posedge 0.1
`define FDM4HSP_SD_PWL 0.1
`define FDM4HSP_CP_PWH 0.1
`define FDM4HSP_CP_PWL 0.1
`define FDM4HSP_D_CP_SETUP_posedge_posedge 0.1
`define FDM4HSP_D_CP_SETUP_negedge_posedge 0.1
`define FDM4HSP_D_CP_HOLD_posedge_posedge 0.1
`define FDM4HSP_D_CP_HOLD_negedge_posedge 0.1

module FDM4HSP (Q, QN, D, CP, SD);

   output Q;
   output QN;
   input D;
   input CP;
   input SD;


   reg Notifier;


   U_FD_P_SN_NOTI u0 (   // Verilog Seq UDP
      IQ, D, CP, SD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   not  (D_, D);

   specify
`ifdef verifault

      if(SD) (posedge CP => (Q +: D)) = (`FDM4HSP_CP_R_Q_R, `FDM4HSP_CP_R_Q_F);
      if(SD) (posedge CP => (QN -: D)) = (`FDM4HSP_CP_R_QN_R, `FDM4HSP_CP_R_QN_F);
      (negedge SD => (Q +: 1'b1)) = (`FDM4HSP_SD_F_Q_R,`FDM4HSP_SD_F_Q_R);
      (negedge SD => (QN +: 1'b0)) = (`FDM4HSP_SD_F_QN_F,`FDM4HSP_SD_F_QN_F);

	$setuphold(posedge CP &&& SD, posedge D, `FDM4HSP_D_CP_SETUP_posedge_posedge, `FDM4HSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& SD, negedge D, `FDM4HSP_D_CP_SETUP_negedge_posedge, `FDM4HSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDM4HSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FDM4HSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FDM4HSP_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_, `FDM4HSP_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_, posedge SD, `FDM4HSP_SD_CP_REM_posedge_posedge, Notifier);


`else
      (posedge CP => (Q +: D)) = (`FDM4HSP_CP_R_Q_R, `FDM4HSP_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`FDM4HSP_CP_R_QN_R, `FDM4HSP_CP_R_QN_F);
      (negedge SD => (Q +: 1'b1)) = (`FDM4HSP_SD_F_Q_R,`FDM4HSP_SD_F_Q_R);
      (negedge SD => (QN +: 1'b0)) = (`FDM4HSP_SD_F_QN_F,`FDM4HSP_SD_F_QN_F);
 
        $setuphold(posedge CP &&& SD, posedge D, `FDM4HSP_D_CP_SETUP_posedge_posedge, `FDM4HSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& SD, negedge D, `FDM4HSP_D_CP_SETUP_negedge_posedge, `FDM4HSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDM4HSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FDM4HSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FDM4HSP_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_, `FDM4HSP_SD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D_, posedge SD, `FDM4HSP_SD_CP_REM_posedge_posedge, Notifier);
 
`endif
   endspecify
`endif


endmodule // FDM4HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:17 and Version :1.1 //
 
//  START 
// CELL FD4QHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD4QHS_SD_F_Q_R 0.1
`define FD4QHS_CP_R_Q_R 0.1
`define FD4QHS_CP_R_Q_F 0.1
`define FD4QHS_D_CP_HOLD_posedge_posedge 0.1
`define FD4QHS_D_CP_HOLD_negedge_posedge 0.1
`define FD4QHS_D_CP_SETUP_posedge_posedge 0.1
`define FD4QHS_D_CP_SETUP_negedge_posedge 0.1
`define FD4QHS_CP_PWL 0.1
`define FD4QHS_CP_PWH 0.1
`define FD4QHS_SD_PWL 0.1
`define FD4QHS_SD_CP_REC_posedge_posedge 0.1
`define FD4QHS_SD_CP_REM_posedge_posedge 0.1

module FD4QHS (Q, D, CP, SD);

   output Q;
   input D;
   input CP;
   input SD;


   reg Notifier;


   U_FD_P_SN_NOTI u0 (IQ, D, CP, SD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   not  (D_, D);

   specify
`ifdef verifault 
      if(SD) (posedge CP => (Q +: D)) = (`FD4QHS_CP_R_Q_R, `FD4QHS_CP_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4QHS_SD_F_Q_R,`FD4QHS_SD_F_Q_R);

	$setuphold(posedge CP &&& SD, posedge D, `FD4QHS_D_CP_SETUP_posedge_posedge, `FD4QHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& SD, negedge D, `FD4QHS_D_CP_SETUP_negedge_posedge, `FD4QHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD4QHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4QHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4QHS_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_, `FD4QHS_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_, posedge SD, `FD4QHS_SD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: D)) = (`FD4QHS_CP_R_Q_R, `FD4QHS_CP_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4QHS_SD_F_Q_R,`FD4QHS_SD_F_Q_R);
 
        $setuphold(posedge CP &&& SD, posedge D, `FD4QHS_D_CP_SETUP_posedge_posedge, `FD4QHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& SD, negedge D, `FD4QHS_D_CP_SETUP_negedge_posedge, `FD4QHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD4QHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4QHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4QHS_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_, `FD4QHS_SD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D_, posedge SD, `FD4QHS_SD_CP_REM_posedge_posedge, Notifier);
 
`endif
   endspecify
`endif


endmodule // FD4QHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:23 and Version :1.1 //
 
//  START 
// CELL FD4QHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD4QHSP_SD_F_Q_R 0.1
`define FD4QHSP_CP_R_Q_R 0.1
`define FD4QHSP_CP_R_Q_F 0.1
`define FD4QHSP_D_CP_HOLD_posedge_posedge 0.1
`define FD4QHSP_D_CP_HOLD_negedge_posedge 0.1
`define FD4QHSP_D_CP_SETUP_posedge_posedge 0.1
`define FD4QHSP_D_CP_SETUP_negedge_posedge 0.1
`define FD4QHSP_CP_PWL 0.1
`define FD4QHSP_CP_PWH 0.1
`define FD4QHSP_SD_PWL 0.1
`define FD4QHSP_SD_CP_REC_posedge_posedge 0.1
`define FD4QHSP_SD_CP_REM_posedge_posedge 0.1

module FD4QHSP (Q, D, CP, SD);

   output Q;
   input D;
   input CP;
   input SD;


   reg Notifier;


   U_FD_P_SN_NOTI u0 (IQ, D, CP, SD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   not  (D_, D);

   specify
`ifdef verifault 
      if(SD) (posedge CP => (Q +: D)) = (`FD4QHSP_CP_R_Q_R, `FD4QHSP_CP_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4QHSP_SD_F_Q_R,`FD4QHSP_SD_F_Q_R);

	$setuphold(posedge CP &&& SD, posedge D, `FD4QHSP_D_CP_SETUP_posedge_posedge, `FD4QHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& SD, negedge D, `FD4QHSP_D_CP_SETUP_negedge_posedge, `FD4QHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD4QHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4QHSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4QHSP_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_, `FD4QHSP_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_, posedge SD, `FD4QHSP_SD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: D)) = (`FD4QHSP_CP_R_Q_R, `FD4QHSP_CP_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4QHSP_SD_F_Q_R,`FD4QHSP_SD_F_Q_R);
 
        $setuphold(posedge CP &&& SD, posedge D, `FD4QHSP_D_CP_SETUP_posedge_posedge, `FD4QHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& SD, negedge D, `FD4QHSP_D_CP_SETUP_negedge_posedge, `FD4QHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD4QHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4QHSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4QHSP_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_, `FD4QHSP_SD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D_, posedge SD, `FD4QHSP_SD_CP_REM_posedge_posedge, Notifier);
 
`endif
   endspecify
`endif


endmodule // FD4QHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:23 and Version :1.1 //
 
//  START 
// CELL FD4QHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD4QHSX4_SD_F_Q_R 0.1
`define FD4QHSX4_CP_R_Q_R 0.1
`define FD4QHSX4_CP_R_Q_F 0.1
`define FD4QHSX4_D_CP_HOLD_posedge_posedge 0.1
`define FD4QHSX4_D_CP_HOLD_negedge_posedge 0.1
`define FD4QHSX4_D_CP_SETUP_posedge_posedge 0.1
`define FD4QHSX4_D_CP_SETUP_negedge_posedge 0.1
`define FD4QHSX4_CP_PWL 0.1
`define FD4QHSX4_CP_PWH 0.1
`define FD4QHSX4_SD_PWL 0.1
`define FD4QHSX4_SD_CP_REC_posedge_posedge 0.1
`define FD4QHSX4_SD_CP_REM_posedge_posedge 0.1

module FD4QHSX4 (Q, D, CP, SD);

   output Q;
   input D;
   input CP;
   input SD;


   reg Notifier;


   U_FD_P_SN_NOTI u0 (IQ, D, CP, SD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   not  (D_, D);

   specify
`ifdef verifault 
      if(SD) (posedge CP => (Q +: D)) = (`FD4QHSX4_CP_R_Q_R, `FD4QHSX4_CP_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4QHSX4_SD_F_Q_R,`FD4QHSX4_SD_F_Q_R);

	$setuphold(posedge CP &&& SD, posedge D, `FD4QHSX4_D_CP_SETUP_posedge_posedge, `FD4QHSX4_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& SD, negedge D, `FD4QHSX4_D_CP_SETUP_negedge_posedge, `FD4QHSX4_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD4QHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4QHSX4_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4QHSX4_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_, `FD4QHSX4_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_, posedge SD, `FD4QHSX4_SD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: D)) = (`FD4QHSX4_CP_R_Q_R, `FD4QHSX4_CP_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4QHSX4_SD_F_Q_R,`FD4QHSX4_SD_F_Q_R);
 
        $setuphold(posedge CP &&& SD, posedge D, `FD4QHSX4_D_CP_SETUP_posedge_posedge, `FD4QHSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& SD, negedge D, `FD4QHSX4_D_CP_SETUP_negedge_posedge, `FD4QHSX4_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD4QHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4QHSX4_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4QHSX4_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_, `FD4QHSX4_SD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D_, posedge SD, `FD4QHSX4_SD_CP_REM_posedge_posedge, Notifier);
 
`endif
   endspecify
`endif


endmodule // FD4QHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:23 and Version :1.1 //
 
//  START 
// CELL FDM4QHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDM4QHS_SD_F_Q_R 0.1
`define FDM4QHS_CP_R_Q_R 0.1
`define FDM4QHS_CP_R_Q_F 0.1
`define FDM4QHS_D_CP_HOLD_posedge_posedge 0.1
`define FDM4QHS_D_CP_HOLD_negedge_posedge 0.1
`define FDM4QHS_D_CP_SETUP_posedge_posedge 0.1
`define FDM4QHS_D_CP_SETUP_negedge_posedge 0.1
`define FDM4QHS_CP_PWL 0.1
`define FDM4QHS_CP_PWH 0.1
`define FDM4QHS_SD_PWL 0.1
`define FDM4QHS_SD_CP_REC_posedge_posedge 0.1
`define FDM4QHS_SD_CP_REM_posedge_posedge 0.1

module FDM4QHS (Q, D, CP, SD);

   output Q;
   input D;
   input CP;
   input SD;


   reg Notifier;


   U_FD_P_SN_NOTI u0 (IQ, D, CP, SD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   not  (D_, D);

   specify
`ifdef verifault 
      if(SD) (posedge CP => (Q +: D)) = (`FDM4QHS_CP_R_Q_R, `FDM4QHS_CP_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FDM4QHS_SD_F_Q_R,`FDM4QHS_SD_F_Q_R);

	$setuphold(posedge CP &&& SD, posedge D, `FDM4QHS_D_CP_SETUP_posedge_posedge, `FDM4QHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& SD, negedge D, `FDM4QHS_D_CP_SETUP_negedge_posedge, `FDM4QHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDM4QHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FDM4QHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FDM4QHS_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_, `FDM4QHS_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_, posedge SD, `FDM4QHS_SD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: D)) = (`FDM4QHS_CP_R_Q_R, `FDM4QHS_CP_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FDM4QHS_SD_F_Q_R,`FDM4QHS_SD_F_Q_R);
 
        $setuphold(posedge CP &&& SD, posedge D, `FDM4QHS_D_CP_SETUP_posedge_posedge, `FDM4QHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& SD, negedge D, `FDM4QHS_D_CP_SETUP_negedge_posedge, `FDM4QHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDM4QHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FDM4QHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FDM4QHS_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_, `FDM4QHS_SD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D_, posedge SD, `FDM4QHS_SD_CP_REM_posedge_posedge, Notifier);
 
`endif
   endspecify
`endif


endmodule // FDM4QHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:23 and Version :1.1 //
 
//  START 
// CELL FDM4QHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDM4QHSP_SD_F_Q_R 0.1
`define FDM4QHSP_CP_R_Q_R 0.1
`define FDM4QHSP_CP_R_Q_F 0.1
`define FDM4QHSP_D_CP_HOLD_posedge_posedge 0.1
`define FDM4QHSP_D_CP_HOLD_negedge_posedge 0.1
`define FDM4QHSP_D_CP_SETUP_posedge_posedge 0.1
`define FDM4QHSP_D_CP_SETUP_negedge_posedge 0.1
`define FDM4QHSP_CP_PWL 0.1
`define FDM4QHSP_CP_PWH 0.1
`define FDM4QHSP_SD_PWL 0.1
`define FDM4QHSP_SD_CP_REC_posedge_posedge 0.1
`define FDM4QHSP_SD_CP_REM_posedge_posedge 0.1

module FDM4QHSP (Q, D, CP, SD);

   output Q;
   input D;
   input CP;
   input SD;


   reg Notifier;


   U_FD_P_SN_NOTI u0 (IQ, D, CP, SD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   not  (D_, D);

   specify
`ifdef verifault 
      if(SD) (posedge CP => (Q +: D)) = (`FDM4QHSP_CP_R_Q_R, `FDM4QHSP_CP_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FDM4QHSP_SD_F_Q_R,`FDM4QHSP_SD_F_Q_R);

	$setuphold(posedge CP &&& SD, posedge D, `FDM4QHSP_D_CP_SETUP_posedge_posedge, `FDM4QHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& SD, negedge D, `FDM4QHSP_D_CP_SETUP_negedge_posedge, `FDM4QHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDM4QHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FDM4QHSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FDM4QHSP_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_, `FDM4QHSP_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_, posedge SD, `FDM4QHSP_SD_CP_REM_posedge_posedge, Notifier);

`else
      (posedge CP => (Q +: D)) = (`FDM4QHSP_CP_R_Q_R, `FDM4QHSP_CP_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FDM4QHSP_SD_F_Q_R,`FDM4QHSP_SD_F_Q_R);
 
        $setuphold(posedge CP &&& SD, posedge D, `FDM4QHSP_D_CP_SETUP_posedge_posedge, `FDM4QHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& SD, negedge D, `FDM4QHSP_D_CP_SETUP_negedge_posedge, `FDM4QHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDM4QHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FDM4QHSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FDM4QHSP_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_, `FDM4QHSP_SD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D_, posedge SD, `FDM4QHSP_SD_CP_REM_posedge_posedge, Notifier);
 
`endif
   endspecify
`endif


endmodule // FDM4QHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:23 and Version :1.1 //
 
//  START 
// CELL FD4SHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD4SHS_SD_F_QN_F 0.1
`define FD4SHS_CP_R_QN_F 0.1
`define FD4SHS_CP_R_QN_R 0.1
`define FD4SHS_SD_F_Q_R 0.1
`define FD4SHS_CP_R_Q_R 0.1
`define FD4SHS_CP_R_Q_F 0.1
`define FD4SHS_SD_CP_REM_posedge_posedge 0.1
`define FD4SHS_SD_CP_REC_posedge_posedge 0.1
`define FD4SHS_SD_PWL 0.1
`define FD4SHS_CP_PWH 0.1
`define FD4SHS_CP_PWL 0.1
`define FD4SHS_D_CP_SETUP_posedge_posedge 0.1
`define FD4SHS_D_CP_SETUP_negedge_posedge 0.1
`define FD4SHS_D_CP_HOLD_posedge_posedge 0.1
`define FD4SHS_D_CP_HOLD_negedge_posedge 0.1
`define FD4SHS_TI_CP_SETUP_posedge_posedge 0.1
`define FD4SHS_TI_CP_SETUP_negedge_posedge 0.1
`define FD4SHS_TI_CP_HOLD_posedge_posedge 0.1
`define FD4SHS_TI_CP_HOLD_negedge_posedge 0.1
`define FD4SHS_TE_CP_SETUP_posedge_posedge 0.1
`define FD4SHS_TE_CP_SETUP_negedge_posedge 0.1
`define FD4SHS_TE_CP_HOLD_posedge_posedge 0.1
`define FD4SHS_TE_CP_HOLD_negedge_posedge 0.1

module FD4SHS (Q, QN, D, CP, SD, TI, TE);

   output Q;
   output QN;
   input D;
   input CP;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_SN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, SD, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   and  (AndSDTEX_, SD, TEX);
   and  (AndSDTE_, SD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_SD_, XorDTI_, SD);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   nor  (D_orTI_onTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && SD) (posedge CP => (Q +: D)) = (`FD4SHS_CP_R_Q_R, `FD4SHS_CP_R_Q_F);
      if(TE && SD) (posedge CP => (Q +: TI)) = (`FD4SHS_CP_R_Q_R, `FD4SHS_CP_R_Q_F);
      if(!D && TI && SD) (posedge CP => (Q +: TE)) = (`FD4SHS_CP_R_Q_R, `FD4SHS_CP_R_Q_F);
      if(!TI && D && SD) (posedge CP => (Q -: TE)) = (`FD4SHS_CP_R_Q_R, `FD4SHS_CP_R_Q_F);
      if(!TE && SD) (posedge CP => (QN -: D)) = (`FD4SHS_CP_R_QN_R, `FD4SHS_CP_R_QN_F);
      if(TE && SD) (posedge CP => (QN -: TI)) = (`FD4SHS_CP_R_QN_R, `FD4SHS_CP_R_QN_F);
      if(!D && TI && SD) (posedge CP => (QN -: TE)) = (`FD4SHS_CP_R_QN_R, `FD4SHS_CP_R_QN_F);
      if(!TI && D && SD) (posedge CP => (QN +: TE)) = (`FD4SHS_CP_R_QN_R, `FD4SHS_CP_R_QN_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4SHS_SD_F_Q_R,`FD4SHS_SD_F_Q_R);
      (negedge SD => (QN +: 1'b0)) = (`FD4SHS_SD_F_QN_F,`FD4SHS_SD_F_QN_F);

	$setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FD4SHS_TE_CP_SETUP_posedge_posedge, `FD4SHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FD4SHS_TE_CP_SETUP_negedge_posedge, `FD4SHS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTE_, posedge TI, `FD4SHS_TI_CP_SETUP_posedge_posedge, `FD4SHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTE_, negedge TI, `FD4SHS_TI_CP_SETUP_negedge_posedge, `FD4SHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTEX_, posedge D, `FD4SHS_D_CP_SETUP_posedge_posedge, `FD4SHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTEX_, negedge D, `FD4SHS_D_CP_SETUP_negedge_posedge, `FD4SHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD4SHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4SHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4SHS_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FD4SHS_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_orTI_onTE, posedge SD, `FD4SHS_SD_CP_REM_posedge_posedge, Notifier);
`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FD4SHS_CP_R_Q_R, `FD4SHS_CP_R_Q_F);
      (posedge CP => (QN -: Mux21DTITE_)) = (`FD4SHS_CP_R_QN_R, `FD4SHS_CP_R_QN_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4SHS_SD_F_Q_R,`FD4SHS_SD_F_Q_R);
      (negedge SD => (QN +: 1'b0)) = (`FD4SHS_SD_F_QN_F,`FD4SHS_SD_F_QN_F);
 
        $setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FD4SHS_TE_CP_SETUP_posedge_posedge, `FD4SHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FD4SHS_TE_CP_SETUP_negedge_posedge, `FD4SHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTE_, posedge TI, `FD4SHS_TI_CP_SETUP_posedge_posedge,`FD4SHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTE_, negedge TI, `FD4SHS_TI_CP_SETUP_negedge_posedge,`FD4SHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTEX_, posedge D, `FD4SHS_D_CP_SETUP_posedge_posedge,`FD4SHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTEX_, negedge D, `FD4SHS_D_CP_SETUP_negedge_posedge,`FD4SHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD4SHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4SHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4SHS_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FD4SHS_SD_CP_REC_posedge_posedge,Notifier);
 
        $hold(posedge CP &&& D_orTI_onTE, posedge SD, `FD4SHS_SD_CP_REM_posedge_posedge, Notifier);

`endif
   endspecify
`endif


endmodule // FD4SHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:27 and Version :1.1 //
 
//  START 
// CELL FD4SHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD4SHSP_SD_F_QN_F 0.1
`define FD4SHSP_CP_R_QN_F 0.1
`define FD4SHSP_CP_R_QN_R 0.1
`define FD4SHSP_SD_F_Q_R 0.1
`define FD4SHSP_CP_R_Q_R 0.1
`define FD4SHSP_CP_R_Q_F 0.1
`define FD4SHSP_SD_CP_REM_posedge_posedge 0.1
`define FD4SHSP_SD_CP_REC_posedge_posedge 0.1
`define FD4SHSP_SD_PWL 0.1
`define FD4SHSP_CP_PWH 0.1
`define FD4SHSP_CP_PWL 0.1
`define FD4SHSP_D_CP_SETUP_posedge_posedge 0.1
`define FD4SHSP_D_CP_SETUP_negedge_posedge 0.1
`define FD4SHSP_D_CP_HOLD_posedge_posedge 0.1
`define FD4SHSP_D_CP_HOLD_negedge_posedge 0.1
`define FD4SHSP_TI_CP_SETUP_posedge_posedge 0.1
`define FD4SHSP_TI_CP_SETUP_negedge_posedge 0.1
`define FD4SHSP_TI_CP_HOLD_posedge_posedge 0.1
`define FD4SHSP_TI_CP_HOLD_negedge_posedge 0.1
`define FD4SHSP_TE_CP_SETUP_posedge_posedge 0.1
`define FD4SHSP_TE_CP_SETUP_negedge_posedge 0.1
`define FD4SHSP_TE_CP_HOLD_posedge_posedge 0.1
`define FD4SHSP_TE_CP_HOLD_negedge_posedge 0.1

module FD4SHSP (Q, QN, D, CP, SD, TI, TE);

   output Q;
   output QN;
   input D;
   input CP;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_SN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, SD, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   and  (AndSDTEX_, SD, TEX);
   and  (AndSDTE_, SD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_SD_, XorDTI_, SD);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   nor  (D_orTI_onTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && SD) (posedge CP => (Q +: D)) = (`FD4SHSP_CP_R_Q_R, `FD4SHSP_CP_R_Q_F);
      if(TE && SD) (posedge CP => (Q +: TI)) = (`FD4SHSP_CP_R_Q_R, `FD4SHSP_CP_R_Q_F);
      if(!D && TI && SD) (posedge CP => (Q +: TE)) = (`FD4SHSP_CP_R_Q_R, `FD4SHSP_CP_R_Q_F);
      if(!TI && D && SD) (posedge CP => (Q -: TE)) = (`FD4SHSP_CP_R_Q_R, `FD4SHSP_CP_R_Q_F);
      if(!TE && SD) (posedge CP => (QN -: D)) = (`FD4SHSP_CP_R_QN_R, `FD4SHSP_CP_R_QN_F);
      if(TE && SD) (posedge CP => (QN -: TI)) = (`FD4SHSP_CP_R_QN_R, `FD4SHSP_CP_R_QN_F);
      if(!D && TI && SD) (posedge CP => (QN -: TE)) = (`FD4SHSP_CP_R_QN_R, `FD4SHSP_CP_R_QN_F);
      if(!TI && D && SD) (posedge CP => (QN +: TE)) = (`FD4SHSP_CP_R_QN_R, `FD4SHSP_CP_R_QN_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4SHSP_SD_F_Q_R,`FD4SHSP_SD_F_Q_R);
      (negedge SD => (QN +: 1'b0)) = (`FD4SHSP_SD_F_QN_F,`FD4SHSP_SD_F_QN_F);

	$setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FD4SHSP_TE_CP_SETUP_posedge_posedge, `FD4SHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FD4SHSP_TE_CP_SETUP_negedge_posedge, `FD4SHSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTE_, posedge TI, `FD4SHSP_TI_CP_SETUP_posedge_posedge, `FD4SHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTE_, negedge TI, `FD4SHSP_TI_CP_SETUP_negedge_posedge, `FD4SHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTEX_, posedge D, `FD4SHSP_D_CP_SETUP_posedge_posedge, `FD4SHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTEX_, negedge D, `FD4SHSP_D_CP_SETUP_negedge_posedge, `FD4SHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD4SHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4SHSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4SHSP_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FD4SHSP_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_orTI_onTE, posedge SD, `FD4SHSP_SD_CP_REM_posedge_posedge, Notifier);
`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FD4SHSP_CP_R_Q_R, `FD4SHSP_CP_R_Q_F);
      (posedge CP => (QN -: Mux21DTITE_)) = (`FD4SHSP_CP_R_QN_R, `FD4SHSP_CP_R_QN_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4SHSP_SD_F_Q_R,`FD4SHSP_SD_F_Q_R);
      (negedge SD => (QN +: 1'b0)) = (`FD4SHSP_SD_F_QN_F,`FD4SHSP_SD_F_QN_F);
 
        $setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FD4SHSP_TE_CP_SETUP_posedge_posedge, `FD4SHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FD4SHSP_TE_CP_SETUP_negedge_posedge, `FD4SHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTE_, posedge TI, `FD4SHSP_TI_CP_SETUP_posedge_posedge,`FD4SHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTE_, negedge TI, `FD4SHSP_TI_CP_SETUP_negedge_posedge,`FD4SHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTEX_, posedge D, `FD4SHSP_D_CP_SETUP_posedge_posedge,`FD4SHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTEX_, negedge D, `FD4SHSP_D_CP_SETUP_negedge_posedge,`FD4SHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD4SHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4SHSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4SHSP_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FD4SHSP_SD_CP_REC_posedge_posedge,Notifier);
 
        $hold(posedge CP &&& D_orTI_onTE, posedge SD, `FD4SHSP_SD_CP_REM_posedge_posedge, Notifier);

`endif
   endspecify
`endif


endmodule // FD4SHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:27 and Version :1.1 //
 
//  START 
// CELL FDM4SHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDM4SHS_SD_F_QN_F 0.1
`define FDM4SHS_CP_R_QN_F 0.1
`define FDM4SHS_CP_R_QN_R 0.1
`define FDM4SHS_SD_F_Q_R 0.1
`define FDM4SHS_CP_R_Q_R 0.1
`define FDM4SHS_CP_R_Q_F 0.1
`define FDM4SHS_SD_CP_REM_posedge_posedge 0.1
`define FDM4SHS_SD_CP_REC_posedge_posedge 0.1
`define FDM4SHS_SD_PWL 0.1
`define FDM4SHS_CP_PWH 0.1
`define FDM4SHS_CP_PWL 0.1
`define FDM4SHS_D_CP_SETUP_posedge_posedge 0.1
`define FDM4SHS_D_CP_SETUP_negedge_posedge 0.1
`define FDM4SHS_D_CP_HOLD_posedge_posedge 0.1
`define FDM4SHS_D_CP_HOLD_negedge_posedge 0.1
`define FDM4SHS_TI_CP_SETUP_posedge_posedge 0.1
`define FDM4SHS_TI_CP_SETUP_negedge_posedge 0.1
`define FDM4SHS_TI_CP_HOLD_posedge_posedge 0.1
`define FDM4SHS_TI_CP_HOLD_negedge_posedge 0.1
`define FDM4SHS_TE_CP_SETUP_posedge_posedge 0.1
`define FDM4SHS_TE_CP_SETUP_negedge_posedge 0.1
`define FDM4SHS_TE_CP_HOLD_posedge_posedge 0.1
`define FDM4SHS_TE_CP_HOLD_negedge_posedge 0.1

module FDM4SHS (Q, QN, D, CP, SD, TI, TE);

   output Q;
   output QN;
   input D;
   input CP;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_SN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, SD, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   and  (AndSDTEX_, SD, TEX);
   and  (AndSDTE_, SD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_SD_, XorDTI_, SD);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   nor  (D_orTI_onTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && SD) (posedge CP => (Q +: D)) = (`FDM4SHS_CP_R_Q_R, `FDM4SHS_CP_R_Q_F);
      if(TE && SD) (posedge CP => (Q +: TI)) = (`FDM4SHS_CP_R_Q_R, `FDM4SHS_CP_R_Q_F);
      if(!D && TI && SD) (posedge CP => (Q +: TE)) = (`FDM4SHS_CP_R_Q_R, `FDM4SHS_CP_R_Q_F);
      if(!TI && D && SD) (posedge CP => (Q -: TE)) = (`FDM4SHS_CP_R_Q_R, `FDM4SHS_CP_R_Q_F);
      if(!TE && SD) (posedge CP => (QN -: D)) = (`FDM4SHS_CP_R_QN_R, `FDM4SHS_CP_R_QN_F);
      if(TE && SD) (posedge CP => (QN -: TI)) = (`FDM4SHS_CP_R_QN_R, `FDM4SHS_CP_R_QN_F);
      if(!D && TI && SD) (posedge CP => (QN -: TE)) = (`FDM4SHS_CP_R_QN_R, `FDM4SHS_CP_R_QN_F);
      if(!TI && D && SD) (posedge CP => (QN +: TE)) = (`FDM4SHS_CP_R_QN_R, `FDM4SHS_CP_R_QN_F);
      (negedge SD => (Q +: 1'b1)) = (`FDM4SHS_SD_F_Q_R,`FDM4SHS_SD_F_Q_R);
      (negedge SD => (QN +: 1'b0)) = (`FDM4SHS_SD_F_QN_F,`FDM4SHS_SD_F_QN_F);

	$setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FDM4SHS_TE_CP_SETUP_posedge_posedge, `FDM4SHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FDM4SHS_TE_CP_SETUP_negedge_posedge, `FDM4SHS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTE_, posedge TI, `FDM4SHS_TI_CP_SETUP_posedge_posedge, `FDM4SHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTE_, negedge TI, `FDM4SHS_TI_CP_SETUP_negedge_posedge, `FDM4SHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTEX_, posedge D, `FDM4SHS_D_CP_SETUP_posedge_posedge, `FDM4SHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTEX_, negedge D, `FDM4SHS_D_CP_SETUP_negedge_posedge, `FDM4SHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDM4SHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FDM4SHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FDM4SHS_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FDM4SHS_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_orTI_onTE, posedge SD, `FDM4SHS_SD_CP_REM_posedge_posedge, Notifier);
`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FDM4SHS_CP_R_Q_R, `FDM4SHS_CP_R_Q_F);
      (posedge CP => (QN -: Mux21DTITE_)) = (`FDM4SHS_CP_R_QN_R, `FDM4SHS_CP_R_QN_F);
      (negedge SD => (Q +: 1'b1)) = (`FDM4SHS_SD_F_Q_R,`FDM4SHS_SD_F_Q_R);
      (negedge SD => (QN +: 1'b0)) = (`FDM4SHS_SD_F_QN_F,`FDM4SHS_SD_F_QN_F);
 
        $setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FDM4SHS_TE_CP_SETUP_posedge_posedge, `FDM4SHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FDM4SHS_TE_CP_SETUP_negedge_posedge, `FDM4SHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTE_, posedge TI, `FDM4SHS_TI_CP_SETUP_posedge_posedge,`FDM4SHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTE_, negedge TI, `FDM4SHS_TI_CP_SETUP_negedge_posedge,`FDM4SHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTEX_, posedge D, `FDM4SHS_D_CP_SETUP_posedge_posedge,`FDM4SHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTEX_, negedge D, `FDM4SHS_D_CP_SETUP_negedge_posedge,`FDM4SHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDM4SHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FDM4SHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FDM4SHS_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FDM4SHS_SD_CP_REC_posedge_posedge,Notifier);
 
        $hold(posedge CP &&& D_orTI_onTE, posedge SD, `FDM4SHS_SD_CP_REM_posedge_posedge, Notifier);

`endif
   endspecify
`endif


endmodule // FDM4SHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:27 and Version :1.1 //
 
//  START 
// CELL FDM4SHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDM4SHSP_SD_F_QN_F 0.1
`define FDM4SHSP_CP_R_QN_F 0.1
`define FDM4SHSP_CP_R_QN_R 0.1
`define FDM4SHSP_SD_F_Q_R 0.1
`define FDM4SHSP_CP_R_Q_R 0.1
`define FDM4SHSP_CP_R_Q_F 0.1
`define FDM4SHSP_SD_CP_REM_posedge_posedge 0.1
`define FDM4SHSP_SD_CP_REC_posedge_posedge 0.1
`define FDM4SHSP_SD_PWL 0.1
`define FDM4SHSP_CP_PWH 0.1
`define FDM4SHSP_CP_PWL 0.1
`define FDM4SHSP_D_CP_SETUP_posedge_posedge 0.1
`define FDM4SHSP_D_CP_SETUP_negedge_posedge 0.1
`define FDM4SHSP_D_CP_HOLD_posedge_posedge 0.1
`define FDM4SHSP_D_CP_HOLD_negedge_posedge 0.1
`define FDM4SHSP_TI_CP_SETUP_posedge_posedge 0.1
`define FDM4SHSP_TI_CP_SETUP_negedge_posedge 0.1
`define FDM4SHSP_TI_CP_HOLD_posedge_posedge 0.1
`define FDM4SHSP_TI_CP_HOLD_negedge_posedge 0.1
`define FDM4SHSP_TE_CP_SETUP_posedge_posedge 0.1
`define FDM4SHSP_TE_CP_SETUP_negedge_posedge 0.1
`define FDM4SHSP_TE_CP_HOLD_posedge_posedge 0.1
`define FDM4SHSP_TE_CP_HOLD_negedge_posedge 0.1

module FDM4SHSP (Q, QN, D, CP, SD, TI, TE);

   output Q;
   output QN;
   input D;
   input CP;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_SN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, SD, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   and  (AndSDTEX_, SD, TEX);
   and  (AndSDTE_, SD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_SD_, XorDTI_, SD);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   nor  (D_orTI_onTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && SD) (posedge CP => (Q +: D)) = (`FDM4SHSP_CP_R_Q_R, `FDM4SHSP_CP_R_Q_F);
      if(TE && SD) (posedge CP => (Q +: TI)) = (`FDM4SHSP_CP_R_Q_R, `FDM4SHSP_CP_R_Q_F);
      if(!D && TI && SD) (posedge CP => (Q +: TE)) = (`FDM4SHSP_CP_R_Q_R, `FDM4SHSP_CP_R_Q_F);
      if(!TI && D && SD) (posedge CP => (Q -: TE)) = (`FDM4SHSP_CP_R_Q_R, `FDM4SHSP_CP_R_Q_F);
      if(!TE && SD) (posedge CP => (QN -: D)) = (`FDM4SHSP_CP_R_QN_R, `FDM4SHSP_CP_R_QN_F);
      if(TE && SD) (posedge CP => (QN -: TI)) = (`FDM4SHSP_CP_R_QN_R, `FDM4SHSP_CP_R_QN_F);
      if(!D && TI && SD) (posedge CP => (QN -: TE)) = (`FDM4SHSP_CP_R_QN_R, `FDM4SHSP_CP_R_QN_F);
      if(!TI && D && SD) (posedge CP => (QN +: TE)) = (`FDM4SHSP_CP_R_QN_R, `FDM4SHSP_CP_R_QN_F);
      (negedge SD => (Q +: 1'b1)) = (`FDM4SHSP_SD_F_Q_R,`FDM4SHSP_SD_F_Q_R);
      (negedge SD => (QN +: 1'b0)) = (`FDM4SHSP_SD_F_QN_F,`FDM4SHSP_SD_F_QN_F);

	$setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FDM4SHSP_TE_CP_SETUP_posedge_posedge, `FDM4SHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FDM4SHSP_TE_CP_SETUP_negedge_posedge, `FDM4SHSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTE_, posedge TI, `FDM4SHSP_TI_CP_SETUP_posedge_posedge, `FDM4SHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTE_, negedge TI, `FDM4SHSP_TI_CP_SETUP_negedge_posedge, `FDM4SHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTEX_, posedge D, `FDM4SHSP_D_CP_SETUP_posedge_posedge, `FDM4SHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTEX_, negedge D, `FDM4SHSP_D_CP_SETUP_negedge_posedge, `FDM4SHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDM4SHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FDM4SHSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FDM4SHSP_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FDM4SHSP_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_orTI_onTE, posedge SD, `FDM4SHSP_SD_CP_REM_posedge_posedge, Notifier);
`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FDM4SHSP_CP_R_Q_R, `FDM4SHSP_CP_R_Q_F);
      (posedge CP => (QN -: Mux21DTITE_)) = (`FDM4SHSP_CP_R_QN_R, `FDM4SHSP_CP_R_QN_F);
      (negedge SD => (Q +: 1'b1)) = (`FDM4SHSP_SD_F_Q_R,`FDM4SHSP_SD_F_Q_R);
      (negedge SD => (QN +: 1'b0)) = (`FDM4SHSP_SD_F_QN_F,`FDM4SHSP_SD_F_QN_F);
 
        $setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FDM4SHSP_TE_CP_SETUP_posedge_posedge, `FDM4SHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FDM4SHSP_TE_CP_SETUP_negedge_posedge, `FDM4SHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTE_, posedge TI, `FDM4SHSP_TI_CP_SETUP_posedge_posedge,`FDM4SHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTE_, negedge TI, `FDM4SHSP_TI_CP_SETUP_negedge_posedge,`FDM4SHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTEX_, posedge D, `FDM4SHSP_D_CP_SETUP_posedge_posedge,`FDM4SHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTEX_, negedge D, `FDM4SHSP_D_CP_SETUP_negedge_posedge,`FDM4SHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDM4SHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FDM4SHSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FDM4SHSP_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FDM4SHSP_SD_CP_REC_posedge_posedge,Notifier);
 
        $hold(posedge CP &&& D_orTI_onTE, posedge SD, `FDM4SHSP_SD_CP_REM_posedge_posedge, Notifier);

`endif
   endspecify
`endif


endmodule // FDM4SHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:27 and Version :1.1 //
 
//  START 
// CELL FD4SQHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD4SQHS_SD_F_Q_R 0.1
`define FD4SQHS_CP_R_Q_R 0.1
`define FD4SQHS_CP_R_Q_F 0.1
`define FD4SQHS_TE_CP_HOLD_posedge_posedge 0.1
`define FD4SQHS_TE_CP_HOLD_negedge_posedge 0.1
`define FD4SQHS_TE_CP_SETUP_posedge_posedge 0.1
`define FD4SQHS_TE_CP_SETUP_negedge_posedge 0.1
`define FD4SQHS_TI_CP_HOLD_posedge_posedge 0.1
`define FD4SQHS_TI_CP_HOLD_negedge_posedge 0.1
`define FD4SQHS_TI_CP_SETUP_posedge_posedge 0.1
`define FD4SQHS_TI_CP_SETUP_negedge_posedge 0.1
`define FD4SQHS_D_CP_HOLD_posedge_posedge 0.1
`define FD4SQHS_D_CP_HOLD_negedge_posedge 0.1
`define FD4SQHS_D_CP_SETUP_posedge_posedge 0.1
`define FD4SQHS_D_CP_SETUP_negedge_posedge 0.1
`define FD4SQHS_CP_PWL 0.1
`define FD4SQHS_CP_PWH 0.1
`define FD4SQHS_SD_PWL 0.1
`define FD4SQHS_SD_CP_REC_posedge_posedge 0.1
`define FD4SQHS_SD_CP_REM_posedge_posedge 0.1

module FD4SQHS (Q, D, CP, SD, TI, TE);

   output Q;
   input D;
   input CP;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_SN_NOTI u1 (IQ, Mux21DTITE_, CP, SD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   and  (AndSDTEX_, SD, TEX);
   not  (TEX, TE);
   and  (AndSDTE_, SD, TE);
   and  (AndXorDTI_SD_, XorDTI_, SD);
   xor  (XorDTI_, D, TI);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   nor  (D_orTI_onTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && SD) (posedge CP => (Q +: D)) = (`FD4SQHS_CP_R_Q_R, `FD4SQHS_CP_R_Q_F);
      if(TE && SD) (posedge CP => (Q +: TI)) = (`FD4SQHS_CP_R_Q_R, `FD4SQHS_CP_R_Q_F);
      if(!D && TI && SD) (posedge CP => (Q +: TE)) = (`FD4SQHS_CP_R_Q_R, `FD4SQHS_CP_R_Q_F);
      if(!TI && D && SD) (posedge CP => (Q -: TE)) = (`FD4SQHS_CP_R_Q_R, `FD4SQHS_CP_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4SQHS_SD_F_Q_R,`FD4SQHS_SD_F_Q_R);

	$setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FD4SQHS_TE_CP_SETUP_posedge_posedge, `FD4SQHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FD4SQHS_TE_CP_SETUP_negedge_posedge, `FD4SQHS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTE_, posedge TI, `FD4SQHS_TI_CP_SETUP_posedge_posedge, `FD4SQHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTE_, negedge TI, `FD4SQHS_TI_CP_SETUP_negedge_posedge, `FD4SQHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTEX_, posedge D, `FD4SQHS_D_CP_SETUP_posedge_posedge, `FD4SQHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTEX_, negedge D, `FD4SQHS_D_CP_SETUP_negedge_posedge, `FD4SQHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD4SQHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4SQHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4SQHS_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FD4SQHS_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_orTI_onTE, posedge SD, `FD4SQHS_SD_CP_REM_posedge_posedge, Notifier);
`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FD4SQHS_CP_R_Q_R, `FD4SQHS_CP_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4SQHS_SD_F_Q_R,`FD4SQHS_SD_F_Q_R);
 
        $setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FD4SQHS_TE_CP_SETUP_posedge_posedge, `FD4SQHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FD4SQHS_TE_CP_SETUP_negedge_posedge, `FD4SQHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTE_, posedge TI, `FD4SQHS_TI_CP_SETUP_posedge_posedge, `FD4SQHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTE_, negedge TI, `FD4SQHS_TI_CP_SETUP_negedge_posedge, `FD4SQHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTEX_, posedge D, `FD4SQHS_D_CP_SETUP_posedge_posedge,`FD4SQHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTEX_, negedge D, `FD4SQHS_D_CP_SETUP_negedge_posedge,`FD4SQHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD4SQHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4SQHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4SQHS_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FD4SQHS_SD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D_orTI_onTE, posedge SD, `FD4SQHS_SD_CP_REM_posedge_posedge, Notifier);

`endif

   endspecify
`endif


endmodule // FD4SQHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:34 and Version :1.1 //
 
//  START 
// CELL FD4SQHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD4SQHSP_SD_F_Q_R 0.1
`define FD4SQHSP_CP_R_Q_R 0.1
`define FD4SQHSP_CP_R_Q_F 0.1
`define FD4SQHSP_TE_CP_HOLD_posedge_posedge 0.1
`define FD4SQHSP_TE_CP_HOLD_negedge_posedge 0.1
`define FD4SQHSP_TE_CP_SETUP_posedge_posedge 0.1
`define FD4SQHSP_TE_CP_SETUP_negedge_posedge 0.1
`define FD4SQHSP_TI_CP_HOLD_posedge_posedge 0.1
`define FD4SQHSP_TI_CP_HOLD_negedge_posedge 0.1
`define FD4SQHSP_TI_CP_SETUP_posedge_posedge 0.1
`define FD4SQHSP_TI_CP_SETUP_negedge_posedge 0.1
`define FD4SQHSP_D_CP_HOLD_posedge_posedge 0.1
`define FD4SQHSP_D_CP_HOLD_negedge_posedge 0.1
`define FD4SQHSP_D_CP_SETUP_posedge_posedge 0.1
`define FD4SQHSP_D_CP_SETUP_negedge_posedge 0.1
`define FD4SQHSP_CP_PWL 0.1
`define FD4SQHSP_CP_PWH 0.1
`define FD4SQHSP_SD_PWL 0.1
`define FD4SQHSP_SD_CP_REC_posedge_posedge 0.1
`define FD4SQHSP_SD_CP_REM_posedge_posedge 0.1

module FD4SQHSP (Q, D, CP, SD, TI, TE);

   output Q;
   input D;
   input CP;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_SN_NOTI u1 (IQ, Mux21DTITE_, CP, SD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   and  (AndSDTEX_, SD, TEX);
   not  (TEX, TE);
   and  (AndSDTE_, SD, TE);
   and  (AndXorDTI_SD_, XorDTI_, SD);
   xor  (XorDTI_, D, TI);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   nor  (D_orTI_onTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && SD) (posedge CP => (Q +: D)) = (`FD4SQHSP_CP_R_Q_R, `FD4SQHSP_CP_R_Q_F);
      if(TE && SD) (posedge CP => (Q +: TI)) = (`FD4SQHSP_CP_R_Q_R, `FD4SQHSP_CP_R_Q_F);
      if(!D && TI && SD) (posedge CP => (Q +: TE)) = (`FD4SQHSP_CP_R_Q_R, `FD4SQHSP_CP_R_Q_F);
      if(!TI && D && SD) (posedge CP => (Q -: TE)) = (`FD4SQHSP_CP_R_Q_R, `FD4SQHSP_CP_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4SQHSP_SD_F_Q_R,`FD4SQHSP_SD_F_Q_R);

	$setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FD4SQHSP_TE_CP_SETUP_posedge_posedge, `FD4SQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FD4SQHSP_TE_CP_SETUP_negedge_posedge, `FD4SQHSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTE_, posedge TI, `FD4SQHSP_TI_CP_SETUP_posedge_posedge, `FD4SQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTE_, negedge TI, `FD4SQHSP_TI_CP_SETUP_negedge_posedge, `FD4SQHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTEX_, posedge D, `FD4SQHSP_D_CP_SETUP_posedge_posedge, `FD4SQHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTEX_, negedge D, `FD4SQHSP_D_CP_SETUP_negedge_posedge, `FD4SQHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD4SQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4SQHSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4SQHSP_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FD4SQHSP_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_orTI_onTE, posedge SD, `FD4SQHSP_SD_CP_REM_posedge_posedge, Notifier);
`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FD4SQHSP_CP_R_Q_R, `FD4SQHSP_CP_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4SQHSP_SD_F_Q_R,`FD4SQHSP_SD_F_Q_R);
 
        $setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FD4SQHSP_TE_CP_SETUP_posedge_posedge, `FD4SQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FD4SQHSP_TE_CP_SETUP_negedge_posedge, `FD4SQHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTE_, posedge TI, `FD4SQHSP_TI_CP_SETUP_posedge_posedge, `FD4SQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTE_, negedge TI, `FD4SQHSP_TI_CP_SETUP_negedge_posedge, `FD4SQHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTEX_, posedge D, `FD4SQHSP_D_CP_SETUP_posedge_posedge,`FD4SQHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTEX_, negedge D, `FD4SQHSP_D_CP_SETUP_negedge_posedge,`FD4SQHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD4SQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4SQHSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4SQHSP_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FD4SQHSP_SD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D_orTI_onTE, posedge SD, `FD4SQHSP_SD_CP_REM_posedge_posedge, Notifier);

`endif

   endspecify
`endif


endmodule // FD4SQHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:34 and Version :1.1 //
 
//  START 
// CELL FD4SQHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD4SQHSX4_SD_F_Q_R 0.1
`define FD4SQHSX4_CP_R_Q_R 0.1
`define FD4SQHSX4_CP_R_Q_F 0.1
`define FD4SQHSX4_TE_CP_HOLD_posedge_posedge 0.1
`define FD4SQHSX4_TE_CP_HOLD_negedge_posedge 0.1
`define FD4SQHSX4_TE_CP_SETUP_posedge_posedge 0.1
`define FD4SQHSX4_TE_CP_SETUP_negedge_posedge 0.1
`define FD4SQHSX4_TI_CP_HOLD_posedge_posedge 0.1
`define FD4SQHSX4_TI_CP_HOLD_negedge_posedge 0.1
`define FD4SQHSX4_TI_CP_SETUP_posedge_posedge 0.1
`define FD4SQHSX4_TI_CP_SETUP_negedge_posedge 0.1
`define FD4SQHSX4_D_CP_HOLD_posedge_posedge 0.1
`define FD4SQHSX4_D_CP_HOLD_negedge_posedge 0.1
`define FD4SQHSX4_D_CP_SETUP_posedge_posedge 0.1
`define FD4SQHSX4_D_CP_SETUP_negedge_posedge 0.1
`define FD4SQHSX4_CP_PWL 0.1
`define FD4SQHSX4_CP_PWH 0.1
`define FD4SQHSX4_SD_PWL 0.1
`define FD4SQHSX4_SD_CP_REC_posedge_posedge 0.1
`define FD4SQHSX4_SD_CP_REM_posedge_posedge 0.1

module FD4SQHSX4 (Q, D, CP, SD, TI, TE);

   output Q;
   input D;
   input CP;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_SN_NOTI u1 (IQ, Mux21DTITE_, CP, SD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   and  (AndSDTEX_, SD, TEX);
   not  (TEX, TE);
   and  (AndSDTE_, SD, TE);
   and  (AndXorDTI_SD_, XorDTI_, SD);
   xor  (XorDTI_, D, TI);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   nor  (D_orTI_onTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && SD) (posedge CP => (Q +: D)) = (`FD4SQHSX4_CP_R_Q_R, `FD4SQHSX4_CP_R_Q_F);
      if(TE && SD) (posedge CP => (Q +: TI)) = (`FD4SQHSX4_CP_R_Q_R, `FD4SQHSX4_CP_R_Q_F);
      if(!D && TI && SD) (posedge CP => (Q +: TE)) = (`FD4SQHSX4_CP_R_Q_R, `FD4SQHSX4_CP_R_Q_F);
      if(!TI && D && SD) (posedge CP => (Q -: TE)) = (`FD4SQHSX4_CP_R_Q_R, `FD4SQHSX4_CP_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4SQHSX4_SD_F_Q_R,`FD4SQHSX4_SD_F_Q_R);

	$setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FD4SQHSX4_TE_CP_SETUP_posedge_posedge, `FD4SQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FD4SQHSX4_TE_CP_SETUP_negedge_posedge, `FD4SQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTE_, posedge TI, `FD4SQHSX4_TI_CP_SETUP_posedge_posedge, `FD4SQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTE_, negedge TI, `FD4SQHSX4_TI_CP_SETUP_negedge_posedge, `FD4SQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTEX_, posedge D, `FD4SQHSX4_D_CP_SETUP_posedge_posedge, `FD4SQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTEX_, negedge D, `FD4SQHSX4_D_CP_SETUP_negedge_posedge, `FD4SQHSX4_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD4SQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4SQHSX4_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4SQHSX4_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FD4SQHSX4_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_orTI_onTE, posedge SD, `FD4SQHSX4_SD_CP_REM_posedge_posedge, Notifier);
`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FD4SQHSX4_CP_R_Q_R, `FD4SQHSX4_CP_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4SQHSX4_SD_F_Q_R,`FD4SQHSX4_SD_F_Q_R);
 
        $setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FD4SQHSX4_TE_CP_SETUP_posedge_posedge, `FD4SQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FD4SQHSX4_TE_CP_SETUP_negedge_posedge, `FD4SQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTE_, posedge TI, `FD4SQHSX4_TI_CP_SETUP_posedge_posedge, `FD4SQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTE_, negedge TI, `FD4SQHSX4_TI_CP_SETUP_negedge_posedge, `FD4SQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTEX_, posedge D, `FD4SQHSX4_D_CP_SETUP_posedge_posedge,`FD4SQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTEX_, negedge D, `FD4SQHSX4_D_CP_SETUP_negedge_posedge,`FD4SQHSX4_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD4SQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4SQHSX4_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4SQHSX4_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FD4SQHSX4_SD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D_orTI_onTE, posedge SD, `FD4SQHSX4_SD_CP_REM_posedge_posedge, Notifier);

`endif

   endspecify
`endif


endmodule // FD4SQHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:34 and Version :1.1 //
 
//  START 
// CELL FDM4SQHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDM4SQHS_SD_F_Q_R 0.1
`define FDM4SQHS_CP_R_Q_R 0.1
`define FDM4SQHS_CP_R_Q_F 0.1
`define FDM4SQHS_TE_CP_HOLD_posedge_posedge 0.1
`define FDM4SQHS_TE_CP_HOLD_negedge_posedge 0.1
`define FDM4SQHS_TE_CP_SETUP_posedge_posedge 0.1
`define FDM4SQHS_TE_CP_SETUP_negedge_posedge 0.1
`define FDM4SQHS_TI_CP_HOLD_posedge_posedge 0.1
`define FDM4SQHS_TI_CP_HOLD_negedge_posedge 0.1
`define FDM4SQHS_TI_CP_SETUP_posedge_posedge 0.1
`define FDM4SQHS_TI_CP_SETUP_negedge_posedge 0.1
`define FDM4SQHS_D_CP_HOLD_posedge_posedge 0.1
`define FDM4SQHS_D_CP_HOLD_negedge_posedge 0.1
`define FDM4SQHS_D_CP_SETUP_posedge_posedge 0.1
`define FDM4SQHS_D_CP_SETUP_negedge_posedge 0.1
`define FDM4SQHS_CP_PWL 0.1
`define FDM4SQHS_CP_PWH 0.1
`define FDM4SQHS_SD_PWL 0.1
`define FDM4SQHS_SD_CP_REC_posedge_posedge 0.1
`define FDM4SQHS_SD_CP_REM_posedge_posedge 0.1

module FDM4SQHS (Q, D, CP, SD, TI, TE);

   output Q;
   input D;
   input CP;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_SN_NOTI u1 (IQ, Mux21DTITE_, CP, SD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   and  (AndSDTEX_, SD, TEX);
   not  (TEX, TE);
   and  (AndSDTE_, SD, TE);
   and  (AndXorDTI_SD_, XorDTI_, SD);
   xor  (XorDTI_, D, TI);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   nor  (D_orTI_onTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && SD) (posedge CP => (Q +: D)) = (`FDM4SQHS_CP_R_Q_R, `FDM4SQHS_CP_R_Q_F);
      if(TE && SD) (posedge CP => (Q +: TI)) = (`FDM4SQHS_CP_R_Q_R, `FDM4SQHS_CP_R_Q_F);
      if(!D && TI && SD) (posedge CP => (Q +: TE)) = (`FDM4SQHS_CP_R_Q_R, `FDM4SQHS_CP_R_Q_F);
      if(!TI && D && SD) (posedge CP => (Q -: TE)) = (`FDM4SQHS_CP_R_Q_R, `FDM4SQHS_CP_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FDM4SQHS_SD_F_Q_R,`FDM4SQHS_SD_F_Q_R);

	$setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FDM4SQHS_TE_CP_SETUP_posedge_posedge, `FDM4SQHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FDM4SQHS_TE_CP_SETUP_negedge_posedge, `FDM4SQHS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTE_, posedge TI, `FDM4SQHS_TI_CP_SETUP_posedge_posedge, `FDM4SQHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTE_, negedge TI, `FDM4SQHS_TI_CP_SETUP_negedge_posedge, `FDM4SQHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTEX_, posedge D, `FDM4SQHS_D_CP_SETUP_posedge_posedge, `FDM4SQHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTEX_, negedge D, `FDM4SQHS_D_CP_SETUP_negedge_posedge, `FDM4SQHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDM4SQHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FDM4SQHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FDM4SQHS_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FDM4SQHS_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_orTI_onTE, posedge SD, `FDM4SQHS_SD_CP_REM_posedge_posedge, Notifier);
`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FDM4SQHS_CP_R_Q_R, `FDM4SQHS_CP_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FDM4SQHS_SD_F_Q_R,`FDM4SQHS_SD_F_Q_R);
 
        $setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FDM4SQHS_TE_CP_SETUP_posedge_posedge, `FDM4SQHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FDM4SQHS_TE_CP_SETUP_negedge_posedge, `FDM4SQHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTE_, posedge TI, `FDM4SQHS_TI_CP_SETUP_posedge_posedge, `FDM4SQHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTE_, negedge TI, `FDM4SQHS_TI_CP_SETUP_negedge_posedge, `FDM4SQHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTEX_, posedge D, `FDM4SQHS_D_CP_SETUP_posedge_posedge,`FDM4SQHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTEX_, negedge D, `FDM4SQHS_D_CP_SETUP_negedge_posedge,`FDM4SQHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDM4SQHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FDM4SQHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FDM4SQHS_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FDM4SQHS_SD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D_orTI_onTE, posedge SD, `FDM4SQHS_SD_CP_REM_posedge_posedge, Notifier);

`endif

   endspecify
`endif


endmodule // FDM4SQHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:34 and Version :1.1 //
 
//  START 
// CELL FDM4SQHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FDM4SQHSP_SD_F_Q_R 0.1
`define FDM4SQHSP_CP_R_Q_R 0.1
`define FDM4SQHSP_CP_R_Q_F 0.1
`define FDM4SQHSP_TE_CP_HOLD_posedge_posedge 0.1
`define FDM4SQHSP_TE_CP_HOLD_negedge_posedge 0.1
`define FDM4SQHSP_TE_CP_SETUP_posedge_posedge 0.1
`define FDM4SQHSP_TE_CP_SETUP_negedge_posedge 0.1
`define FDM4SQHSP_TI_CP_HOLD_posedge_posedge 0.1
`define FDM4SQHSP_TI_CP_HOLD_negedge_posedge 0.1
`define FDM4SQHSP_TI_CP_SETUP_posedge_posedge 0.1
`define FDM4SQHSP_TI_CP_SETUP_negedge_posedge 0.1
`define FDM4SQHSP_D_CP_HOLD_posedge_posedge 0.1
`define FDM4SQHSP_D_CP_HOLD_negedge_posedge 0.1
`define FDM4SQHSP_D_CP_SETUP_posedge_posedge 0.1
`define FDM4SQHSP_D_CP_SETUP_negedge_posedge 0.1
`define FDM4SQHSP_CP_PWL 0.1
`define FDM4SQHSP_CP_PWH 0.1
`define FDM4SQHSP_SD_PWL 0.1
`define FDM4SQHSP_SD_CP_REC_posedge_posedge 0.1
`define FDM4SQHSP_SD_CP_REM_posedge_posedge 0.1

module FDM4SQHSP (Q, D, CP, SD, TI, TE);

   output Q;
   input D;
   input CP;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_SN_NOTI u1 (IQ, Mux21DTITE_, CP, SD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   and  (AndSDTEX_, SD, TEX);
   not  (TEX, TE);
   and  (AndSDTE_, SD, TE);
   and  (AndXorDTI_SD_, XorDTI_, SD);
   xor  (XorDTI_, D, TI);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   nor  (D_orTI_onTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && SD) (posedge CP => (Q +: D)) = (`FDM4SQHSP_CP_R_Q_R, `FDM4SQHSP_CP_R_Q_F);
      if(TE && SD) (posedge CP => (Q +: TI)) = (`FDM4SQHSP_CP_R_Q_R, `FDM4SQHSP_CP_R_Q_F);
      if(!D && TI && SD) (posedge CP => (Q +: TE)) = (`FDM4SQHSP_CP_R_Q_R, `FDM4SQHSP_CP_R_Q_F);
      if(!TI && D && SD) (posedge CP => (Q -: TE)) = (`FDM4SQHSP_CP_R_Q_R, `FDM4SQHSP_CP_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FDM4SQHSP_SD_F_Q_R,`FDM4SQHSP_SD_F_Q_R);

	$setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FDM4SQHSP_TE_CP_SETUP_posedge_posedge, `FDM4SQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FDM4SQHSP_TE_CP_SETUP_negedge_posedge, `FDM4SQHSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTE_, posedge TI, `FDM4SQHSP_TI_CP_SETUP_posedge_posedge, `FDM4SQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTE_, negedge TI, `FDM4SQHSP_TI_CP_SETUP_negedge_posedge, `FDM4SQHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTEX_, posedge D, `FDM4SQHSP_D_CP_SETUP_posedge_posedge, `FDM4SQHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTEX_, negedge D, `FDM4SQHSP_D_CP_SETUP_negedge_posedge, `FDM4SQHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FDM4SQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FDM4SQHSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FDM4SQHSP_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FDM4SQHSP_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_orTI_onTE, posedge SD, `FDM4SQHSP_SD_CP_REM_posedge_posedge, Notifier);
`else
      (posedge CP => (Q +: Mux21DTITE_)) = (`FDM4SQHSP_CP_R_Q_R, `FDM4SQHSP_CP_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FDM4SQHSP_SD_F_Q_R,`FDM4SQHSP_SD_F_Q_R);
 
        $setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FDM4SQHSP_TE_CP_SETUP_posedge_posedge, `FDM4SQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FDM4SQHSP_TE_CP_SETUP_negedge_posedge, `FDM4SQHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTE_, posedge TI, `FDM4SQHSP_TI_CP_SETUP_posedge_posedge, `FDM4SQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTE_, negedge TI, `FDM4SQHSP_TI_CP_SETUP_negedge_posedge, `FDM4SQHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTEX_, posedge D, `FDM4SQHSP_D_CP_SETUP_posedge_posedge,`FDM4SQHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTEX_, negedge D, `FDM4SQHSP_D_CP_SETUP_negedge_posedge,`FDM4SQHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FDM4SQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FDM4SQHSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FDM4SQHSP_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FDM4SQHSP_SD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D_orTI_onTE, posedge SD, `FDM4SQHSP_SD_CP_REM_posedge_posedge, Notifier);

`endif

   endspecify
`endif


endmodule // FDM4SQHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:34 and Version :1.1 //
 
//  START 
// CELL FD4THS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD4THS_SD_F_SO_R 0.1
`define FD4THS_CP_R_SO_R 0.1
`define FD4THS_CP_R_SO_F 0.1
`define FD4THS_SD_F_QN_F 0.1
`define FD4THS_CP_R_QN_F 0.1
`define FD4THS_CP_R_QN_R 0.1
`define FD4THS_SD_F_Q_R 0.1
`define FD4THS_CP_R_Q_R 0.1
`define FD4THS_CP_R_Q_F 0.1
`define FD4THS_SD_CP_REM_posedge_posedge 0.1
`define FD4THS_SD_CP_REC_posedge_posedge 0.1
`define FD4THS_SD_PWL 0.1
`define FD4THS_CP_PWH 0.1
`define FD4THS_CP_PWL 0.1
`define FD4THS_D_CP_SETUP_posedge_posedge 0.1
`define FD4THS_D_CP_SETUP_negedge_posedge 0.1
`define FD4THS_D_CP_HOLD_posedge_posedge 0.1
`define FD4THS_D_CP_HOLD_negedge_posedge 0.1
`define FD4THS_TI_CP_SETUP_posedge_posedge 0.1
`define FD4THS_TI_CP_SETUP_negedge_posedge 0.1
`define FD4THS_TI_CP_HOLD_posedge_posedge 0.1
`define FD4THS_TI_CP_HOLD_negedge_posedge 0.1
`define FD4THS_TE_CP_SETUP_posedge_posedge 0.1
`define FD4THS_TE_CP_SETUP_negedge_posedge 0.1
`define FD4THS_TE_CP_HOLD_posedge_posedge 0.1
`define FD4THS_TE_CP_HOLD_negedge_posedge 0.1

module FD4THS (Q, QN, SO, D, CP, SD, TI, TE);

   output Q;
   output QN;
   output SO;
   input D;
   input CP;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_SN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, SD, Notifier);

   buf  u2 (Q, IQ);
   buf  u3 (SO, IQ);
   not  u4 (QN, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   and  (AndSDTEX_, SD, TEX);
   and  (AndSDTE_, SD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_SD_, XorDTI_, SD);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   nor  (D_orTI_onTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && SD) (posedge CP => (Q +: D)) = (`FD4THS_CP_R_Q_R, `FD4THS_CP_R_Q_F);
      if(TE && SD) (posedge CP => (Q +: TI)) = (`FD4THS_CP_R_Q_R, `FD4THS_CP_R_Q_F);
      if(!D && TI && SD) (posedge CP => (Q +: TE)) = (`FD4THS_CP_R_Q_R, `FD4THS_CP_R_Q_F);
      if(!TI && D && SD) (posedge CP => (Q -: TE)) = (`FD4THS_CP_R_Q_R, `FD4THS_CP_R_Q_F);
      if(!TE && SD) (posedge CP => (QN -: D)) = (`FD4THS_CP_R_QN_R, `FD4THS_CP_R_QN_F);
      if(TE && SD) (posedge CP => (QN -: TI)) = (`FD4THS_CP_R_QN_R, `FD4THS_CP_R_QN_F);
      if(!D && TI && SD) (posedge CP => (QN -: TE)) = (`FD4THS_CP_R_QN_R, `FD4THS_CP_R_QN_F);
      if(!TI && D && SD) (posedge CP => (QN +: TE)) = (`FD4THS_CP_R_QN_R, `FD4THS_CP_R_QN_F);
      if(!TE && SD) (posedge CP => (SO +: D)) = (`FD4THS_CP_R_SO_R, `FD4THS_CP_R_SO_F);
      if(TE && SD) (posedge CP => (SO +: TI)) = (`FD4THS_CP_R_SO_R, `FD4THS_CP_R_SO_F);
      if(!D && TI && SD) (posedge CP => (SO +: TE)) = (`FD4THS_CP_R_SO_R, `FD4THS_CP_R_SO_F);
      if(!TI && D && SD) (posedge CP => (SO -: TE)) = (`FD4THS_CP_R_SO_R, `FD4THS_CP_R_SO_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4THS_SD_F_Q_R,`FD4THS_SD_F_Q_R);
      (negedge SD => (QN +: 1'b0)) = (`FD4THS_SD_F_QN_F,`FD4THS_SD_F_QN_F);
      (negedge SD => (SO +: 1'b1)) = (`FD4THS_SD_F_SO_R,`FD4THS_SD_F_SO_R);

	$setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FD4THS_TE_CP_SETUP_posedge_posedge, `FD4THS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FD4THS_TE_CP_SETUP_negedge_posedge, `FD4THS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTE_, posedge TI, `FD4THS_TI_CP_SETUP_posedge_posedge, `FD4THS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTE_, negedge TI, `FD4THS_TI_CP_SETUP_negedge_posedge, `FD4THS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTEX_, posedge D, `FD4THS_D_CP_SETUP_posedge_posedge, `FD4THS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTEX_, negedge D, `FD4THS_D_CP_SETUP_negedge_posedge, `FD4THS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD4THS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4THS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4THS_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FD4THS_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_orTI_onTE, posedge SD, `FD4THS_SD_CP_REM_posedge_posedge, Notifier);

`else

      (posedge CP => (Q +: Mux21DTITE_)) = (`FD4THS_CP_R_Q_R, `FD4THS_CP_R_Q_F);
      (posedge CP => (QN -: Mux21DTITE_)) = (`FD4THS_CP_R_QN_R, `FD4THS_CP_R_QN_F);
      (posedge CP => (SO +: Mux21DTITE_)) = (`FD4THS_CP_R_SO_R, `FD4THS_CP_R_SO_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4THS_SD_F_Q_R,`FD4THS_SD_F_Q_R);
      (negedge SD => (QN +: 1'b0)) = (`FD4THS_SD_F_QN_F,`FD4THS_SD_F_QN_F);
      (negedge SD => (SO +: 1'b1)) = (`FD4THS_SD_F_SO_R,`FD4THS_SD_F_SO_R);
 
        $setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FD4THS_TE_CP_SETUP_posedge_posedge, `FD4THS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FD4THS_TE_CP_SETUP_negedge_posedge, `FD4THS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTE_, posedge TI, `FD4THS_TI_CP_SETUP_posedge_posedge, `FD4THS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTE_, negedge TI, `FD4THS_TI_CP_SETUP_negedge_posedge, `FD4THS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTEX_, posedge D, `FD4THS_D_CP_SETUP_posedge_posedge, `FD4THS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTEX_, negedge D, `FD4THS_D_CP_SETUP_negedge_posedge, `FD4THS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD4THS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4THS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4THS_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FD4THS_SD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D_orTI_onTE, posedge SD, `FD4THS_SD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FD4THS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:38 and Version :1.1 //
 
//  START 
// CELL FD4THSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD4THSP_SD_F_SO_R 0.1
`define FD4THSP_CP_R_SO_R 0.1
`define FD4THSP_CP_R_SO_F 0.1
`define FD4THSP_SD_F_QN_F 0.1
`define FD4THSP_CP_R_QN_F 0.1
`define FD4THSP_CP_R_QN_R 0.1
`define FD4THSP_SD_F_Q_R 0.1
`define FD4THSP_CP_R_Q_R 0.1
`define FD4THSP_CP_R_Q_F 0.1
`define FD4THSP_SD_CP_REM_posedge_posedge 0.1
`define FD4THSP_SD_CP_REC_posedge_posedge 0.1
`define FD4THSP_SD_PWL 0.1
`define FD4THSP_CP_PWH 0.1
`define FD4THSP_CP_PWL 0.1
`define FD4THSP_D_CP_SETUP_posedge_posedge 0.1
`define FD4THSP_D_CP_SETUP_negedge_posedge 0.1
`define FD4THSP_D_CP_HOLD_posedge_posedge 0.1
`define FD4THSP_D_CP_HOLD_negedge_posedge 0.1
`define FD4THSP_TI_CP_SETUP_posedge_posedge 0.1
`define FD4THSP_TI_CP_SETUP_negedge_posedge 0.1
`define FD4THSP_TI_CP_HOLD_posedge_posedge 0.1
`define FD4THSP_TI_CP_HOLD_negedge_posedge 0.1
`define FD4THSP_TE_CP_SETUP_posedge_posedge 0.1
`define FD4THSP_TE_CP_SETUP_negedge_posedge 0.1
`define FD4THSP_TE_CP_HOLD_posedge_posedge 0.1
`define FD4THSP_TE_CP_HOLD_negedge_posedge 0.1

module FD4THSP (Q, QN, SO, D, CP, SD, TI, TE);

   output Q;
   output QN;
   output SO;
   input D;
   input CP;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_SN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, SD, Notifier);

   buf  u2 (Q, IQ);
   buf  u3 (SO, IQ);
   not  u4 (QN, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   and  (AndSDTEX_, SD, TEX);
   and  (AndSDTE_, SD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_SD_, XorDTI_, SD);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   nor  (D_orTI_onTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && SD) (posedge CP => (Q +: D)) = (`FD4THSP_CP_R_Q_R, `FD4THSP_CP_R_Q_F);
      if(TE && SD) (posedge CP => (Q +: TI)) = (`FD4THSP_CP_R_Q_R, `FD4THSP_CP_R_Q_F);
      if(!D && TI && SD) (posedge CP => (Q +: TE)) = (`FD4THSP_CP_R_Q_R, `FD4THSP_CP_R_Q_F);
      if(!TI && D && SD) (posedge CP => (Q -: TE)) = (`FD4THSP_CP_R_Q_R, `FD4THSP_CP_R_Q_F);
      if(!TE && SD) (posedge CP => (QN -: D)) = (`FD4THSP_CP_R_QN_R, `FD4THSP_CP_R_QN_F);
      if(TE && SD) (posedge CP => (QN -: TI)) = (`FD4THSP_CP_R_QN_R, `FD4THSP_CP_R_QN_F);
      if(!D && TI && SD) (posedge CP => (QN -: TE)) = (`FD4THSP_CP_R_QN_R, `FD4THSP_CP_R_QN_F);
      if(!TI && D && SD) (posedge CP => (QN +: TE)) = (`FD4THSP_CP_R_QN_R, `FD4THSP_CP_R_QN_F);
      if(!TE && SD) (posedge CP => (SO +: D)) = (`FD4THSP_CP_R_SO_R, `FD4THSP_CP_R_SO_F);
      if(TE && SD) (posedge CP => (SO +: TI)) = (`FD4THSP_CP_R_SO_R, `FD4THSP_CP_R_SO_F);
      if(!D && TI && SD) (posedge CP => (SO +: TE)) = (`FD4THSP_CP_R_SO_R, `FD4THSP_CP_R_SO_F);
      if(!TI && D && SD) (posedge CP => (SO -: TE)) = (`FD4THSP_CP_R_SO_R, `FD4THSP_CP_R_SO_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4THSP_SD_F_Q_R,`FD4THSP_SD_F_Q_R);
      (negedge SD => (QN +: 1'b0)) = (`FD4THSP_SD_F_QN_F,`FD4THSP_SD_F_QN_F);
      (negedge SD => (SO +: 1'b1)) = (`FD4THSP_SD_F_SO_R,`FD4THSP_SD_F_SO_R);

	$setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FD4THSP_TE_CP_SETUP_posedge_posedge, `FD4THSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FD4THSP_TE_CP_SETUP_negedge_posedge, `FD4THSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTE_, posedge TI, `FD4THSP_TI_CP_SETUP_posedge_posedge, `FD4THSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTE_, negedge TI, `FD4THSP_TI_CP_SETUP_negedge_posedge, `FD4THSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTEX_, posedge D, `FD4THSP_D_CP_SETUP_posedge_posedge, `FD4THSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTEX_, negedge D, `FD4THSP_D_CP_SETUP_negedge_posedge, `FD4THSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD4THSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4THSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4THSP_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FD4THSP_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_orTI_onTE, posedge SD, `FD4THSP_SD_CP_REM_posedge_posedge, Notifier);

`else

      (posedge CP => (Q +: Mux21DTITE_)) = (`FD4THSP_CP_R_Q_R, `FD4THSP_CP_R_Q_F);
      (posedge CP => (QN -: Mux21DTITE_)) = (`FD4THSP_CP_R_QN_R, `FD4THSP_CP_R_QN_F);
      (posedge CP => (SO +: Mux21DTITE_)) = (`FD4THSP_CP_R_SO_R, `FD4THSP_CP_R_SO_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4THSP_SD_F_Q_R,`FD4THSP_SD_F_Q_R);
      (negedge SD => (QN +: 1'b0)) = (`FD4THSP_SD_F_QN_F,`FD4THSP_SD_F_QN_F);
      (negedge SD => (SO +: 1'b1)) = (`FD4THSP_SD_F_SO_R,`FD4THSP_SD_F_SO_R);
 
        $setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FD4THSP_TE_CP_SETUP_posedge_posedge, `FD4THSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FD4THSP_TE_CP_SETUP_negedge_posedge, `FD4THSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTE_, posedge TI, `FD4THSP_TI_CP_SETUP_posedge_posedge, `FD4THSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTE_, negedge TI, `FD4THSP_TI_CP_SETUP_negedge_posedge, `FD4THSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTEX_, posedge D, `FD4THSP_D_CP_SETUP_posedge_posedge, `FD4THSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTEX_, negedge D, `FD4THSP_D_CP_SETUP_negedge_posedge, `FD4THSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD4THSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4THSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4THSP_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FD4THSP_SD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D_orTI_onTE, posedge SD, `FD4THSP_SD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FD4THSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:38 and Version :1.1 //
 
//  START 
// CELL FD4TQHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD4TQHS_SD_F_SO_R 0.1
`define FD4TQHS_CP_R_SO_R 0.1
`define FD4TQHS_CP_R_SO_F 0.1
`define FD4TQHS_SD_F_Q_R 0.1
`define FD4TQHS_CP_R_Q_R 0.1
`define FD4TQHS_CP_R_Q_F 0.1
`define FD4TQHS_SD_CP_REM_posedge_posedge 0.1
`define FD4TQHS_SD_CP_REC_posedge_posedge 0.1
`define FD4TQHS_SD_PWL 0.1
`define FD4TQHS_CP_PWH 0.1
`define FD4TQHS_CP_PWL 0.1
`define FD4TQHS_D_CP_SETUP_posedge_posedge 0.1
`define FD4TQHS_D_CP_SETUP_negedge_posedge 0.1
`define FD4TQHS_D_CP_HOLD_posedge_posedge 0.1
`define FD4TQHS_D_CP_HOLD_negedge_posedge 0.1
`define FD4TQHS_TI_CP_SETUP_posedge_posedge 0.1
`define FD4TQHS_TI_CP_SETUP_negedge_posedge 0.1
`define FD4TQHS_TI_CP_HOLD_posedge_posedge 0.1
`define FD4TQHS_TI_CP_HOLD_negedge_posedge 0.1
`define FD4TQHS_TE_CP_SETUP_posedge_posedge 0.1
`define FD4TQHS_TE_CP_SETUP_negedge_posedge 0.1
`define FD4TQHS_TE_CP_HOLD_posedge_posedge 0.1
`define FD4TQHS_TE_CP_HOLD_negedge_posedge 0.1

module FD4TQHS (Q, SO, D, CP, SD, TI, TE);

   output Q;
   output SO;
   input D;
   input CP;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_SN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, SD, Notifier);

   buf  u2 (Q, IQ);
   buf  u3 (SO, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   and  (AndSDTEX_, SD, TEX);
   and  (AndSDTE_, SD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_SD_, XorDTI_, SD);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   nor  (D_orTI_onTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && SD) (posedge CP => (Q +: D)) = (`FD4TQHS_CP_R_Q_R, `FD4TQHS_CP_R_Q_F);
      if(TE && SD) (posedge CP => (Q +: TI)) = (`FD4TQHS_CP_R_Q_R, `FD4TQHS_CP_R_Q_F);
      if(!D && TI && SD) (posedge CP => (Q +: TE)) = (`FD4TQHS_CP_R_Q_R, `FD4TQHS_CP_R_Q_F);
      if(!TI && D && SD) (posedge CP => (Q -: TE)) = (`FD4TQHS_CP_R_Q_R, `FD4TQHS_CP_R_Q_F);
      if(!TE && SD) (posedge CP => (SO +: D)) = (`FD4TQHS_CP_R_SO_R, `FD4TQHS_CP_R_SO_F);
      if(TE && SD) (posedge CP => (SO +: TI)) = (`FD4TQHS_CP_R_SO_R, `FD4TQHS_CP_R_SO_F);
      if(!D && TI && SD) (posedge CP => (SO +: TE)) = (`FD4TQHS_CP_R_SO_R, `FD4TQHS_CP_R_SO_F);
      if(!TI && D && SD) (posedge CP => (SO -: TE)) = (`FD4TQHS_CP_R_SO_R, `FD4TQHS_CP_R_SO_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4TQHS_SD_F_Q_R,`FD4TQHS_SD_F_Q_R);
      (negedge SD => (SO +: 1'b1)) = (`FD4TQHS_SD_F_SO_R,`FD4TQHS_SD_F_SO_R);

	$setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FD4TQHS_TE_CP_SETUP_posedge_posedge, `FD4TQHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FD4TQHS_TE_CP_SETUP_negedge_posedge, `FD4TQHS_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTE_, posedge TI, `FD4TQHS_TI_CP_SETUP_posedge_posedge, `FD4TQHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTE_, negedge TI, `FD4TQHS_TI_CP_SETUP_negedge_posedge, `FD4TQHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTEX_, posedge D, `FD4TQHS_D_CP_SETUP_posedge_posedge, `FD4TQHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTEX_, negedge D, `FD4TQHS_D_CP_SETUP_negedge_posedge, `FD4TQHS_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD4TQHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4TQHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4TQHS_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FD4TQHS_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_orTI_onTE, posedge SD, `FD4TQHS_SD_CP_REM_posedge_posedge, Notifier);
`else
       (posedge CP => (Q +: Mux21DTITE_)) = (`FD4TQHS_CP_R_Q_R, `FD4TQHS_CP_R_Q_F);
       (posedge CP => (SO +: Mux21DTITE_)) = (`FD4TQHS_CP_R_SO_R, `FD4TQHS_CP_R_SO_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4TQHS_SD_F_Q_R,`FD4TQHS_SD_F_Q_R);
      (negedge SD => (SO +: 1'b1)) = (`FD4TQHS_SD_F_SO_R,`FD4TQHS_SD_F_SO_R);
 
        $setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FD4TQHS_TE_CP_SETUP_posedge_posedge, `FD4TQHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FD4TQHS_TE_CP_SETUP_negedge_posedge, `FD4TQHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTE_, posedge TI, `FD4TQHS_TI_CP_SETUP_posedge_posedge, `FD4TQHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTE_, negedge TI, `FD4TQHS_TI_CP_SETUP_negedge_posedge, `FD4TQHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTEX_, posedge D, `FD4TQHS_D_CP_SETUP_posedge_posedge,`FD4TQHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTEX_, negedge D, `FD4TQHS_D_CP_SETUP_negedge_posedge,`FD4TQHS_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD4TQHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4TQHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4TQHS_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FD4TQHS_SD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D_orTI_onTE, posedge SD, `FD4TQHS_SD_CP_REM_posedge_posedge, Notifier);

`endif

   endspecify
`endif


endmodule // FD4TQHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:44 and Version :1.1 //
 
//  START 
// CELL FD4TQHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD4TQHSP_SD_F_SO_R 0.1
`define FD4TQHSP_CP_R_SO_R 0.1
`define FD4TQHSP_CP_R_SO_F 0.1
`define FD4TQHSP_SD_F_Q_R 0.1
`define FD4TQHSP_CP_R_Q_R 0.1
`define FD4TQHSP_CP_R_Q_F 0.1
`define FD4TQHSP_SD_CP_REM_posedge_posedge 0.1
`define FD4TQHSP_SD_CP_REC_posedge_posedge 0.1
`define FD4TQHSP_SD_PWL 0.1
`define FD4TQHSP_CP_PWH 0.1
`define FD4TQHSP_CP_PWL 0.1
`define FD4TQHSP_D_CP_SETUP_posedge_posedge 0.1
`define FD4TQHSP_D_CP_SETUP_negedge_posedge 0.1
`define FD4TQHSP_D_CP_HOLD_posedge_posedge 0.1
`define FD4TQHSP_D_CP_HOLD_negedge_posedge 0.1
`define FD4TQHSP_TI_CP_SETUP_posedge_posedge 0.1
`define FD4TQHSP_TI_CP_SETUP_negedge_posedge 0.1
`define FD4TQHSP_TI_CP_HOLD_posedge_posedge 0.1
`define FD4TQHSP_TI_CP_HOLD_negedge_posedge 0.1
`define FD4TQHSP_TE_CP_SETUP_posedge_posedge 0.1
`define FD4TQHSP_TE_CP_SETUP_negedge_posedge 0.1
`define FD4TQHSP_TE_CP_HOLD_posedge_posedge 0.1
`define FD4TQHSP_TE_CP_HOLD_negedge_posedge 0.1

module FD4TQHSP (Q, SO, D, CP, SD, TI, TE);

   output Q;
   output SO;
   input D;
   input CP;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_SN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, SD, Notifier);

   buf  u2 (Q, IQ);
   buf  u3 (SO, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   and  (AndSDTEX_, SD, TEX);
   and  (AndSDTE_, SD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_SD_, XorDTI_, SD);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   nor  (D_orTI_onTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && SD) (posedge CP => (Q +: D)) = (`FD4TQHSP_CP_R_Q_R, `FD4TQHSP_CP_R_Q_F);
      if(TE && SD) (posedge CP => (Q +: TI)) = (`FD4TQHSP_CP_R_Q_R, `FD4TQHSP_CP_R_Q_F);
      if(!D && TI && SD) (posedge CP => (Q +: TE)) = (`FD4TQHSP_CP_R_Q_R, `FD4TQHSP_CP_R_Q_F);
      if(!TI && D && SD) (posedge CP => (Q -: TE)) = (`FD4TQHSP_CP_R_Q_R, `FD4TQHSP_CP_R_Q_F);
      if(!TE && SD) (posedge CP => (SO +: D)) = (`FD4TQHSP_CP_R_SO_R, `FD4TQHSP_CP_R_SO_F);
      if(TE && SD) (posedge CP => (SO +: TI)) = (`FD4TQHSP_CP_R_SO_R, `FD4TQHSP_CP_R_SO_F);
      if(!D && TI && SD) (posedge CP => (SO +: TE)) = (`FD4TQHSP_CP_R_SO_R, `FD4TQHSP_CP_R_SO_F);
      if(!TI && D && SD) (posedge CP => (SO -: TE)) = (`FD4TQHSP_CP_R_SO_R, `FD4TQHSP_CP_R_SO_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4TQHSP_SD_F_Q_R,`FD4TQHSP_SD_F_Q_R);
      (negedge SD => (SO +: 1'b1)) = (`FD4TQHSP_SD_F_SO_R,`FD4TQHSP_SD_F_SO_R);

	$setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FD4TQHSP_TE_CP_SETUP_posedge_posedge, `FD4TQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FD4TQHSP_TE_CP_SETUP_negedge_posedge, `FD4TQHSP_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTE_, posedge TI, `FD4TQHSP_TI_CP_SETUP_posedge_posedge, `FD4TQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTE_, negedge TI, `FD4TQHSP_TI_CP_SETUP_negedge_posedge, `FD4TQHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTEX_, posedge D, `FD4TQHSP_D_CP_SETUP_posedge_posedge, `FD4TQHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTEX_, negedge D, `FD4TQHSP_D_CP_SETUP_negedge_posedge, `FD4TQHSP_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD4TQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4TQHSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4TQHSP_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FD4TQHSP_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_orTI_onTE, posedge SD, `FD4TQHSP_SD_CP_REM_posedge_posedge, Notifier);
`else
       (posedge CP => (Q +: Mux21DTITE_)) = (`FD4TQHSP_CP_R_Q_R, `FD4TQHSP_CP_R_Q_F);
       (posedge CP => (SO +: Mux21DTITE_)) = (`FD4TQHSP_CP_R_SO_R, `FD4TQHSP_CP_R_SO_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4TQHSP_SD_F_Q_R,`FD4TQHSP_SD_F_Q_R);
      (negedge SD => (SO +: 1'b1)) = (`FD4TQHSP_SD_F_SO_R,`FD4TQHSP_SD_F_SO_R);
 
        $setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FD4TQHSP_TE_CP_SETUP_posedge_posedge, `FD4TQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FD4TQHSP_TE_CP_SETUP_negedge_posedge, `FD4TQHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTE_, posedge TI, `FD4TQHSP_TI_CP_SETUP_posedge_posedge, `FD4TQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTE_, negedge TI, `FD4TQHSP_TI_CP_SETUP_negedge_posedge, `FD4TQHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTEX_, posedge D, `FD4TQHSP_D_CP_SETUP_posedge_posedge,`FD4TQHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTEX_, negedge D, `FD4TQHSP_D_CP_SETUP_negedge_posedge,`FD4TQHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD4TQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4TQHSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4TQHSP_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FD4TQHSP_SD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D_orTI_onTE, posedge SD, `FD4TQHSP_SD_CP_REM_posedge_posedge, Notifier);

`endif

   endspecify
`endif


endmodule // FD4TQHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:44 and Version :1.1 //
 
//  START 
// CELL FD4TQHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD4TQHSX4_SD_F_SO_R 0.1
`define FD4TQHSX4_CP_R_SO_R 0.1
`define FD4TQHSX4_CP_R_SO_F 0.1
`define FD4TQHSX4_SD_F_Q_R 0.1
`define FD4TQHSX4_CP_R_Q_R 0.1
`define FD4TQHSX4_CP_R_Q_F 0.1
`define FD4TQHSX4_SD_CP_REM_posedge_posedge 0.1
`define FD4TQHSX4_SD_CP_REC_posedge_posedge 0.1
`define FD4TQHSX4_SD_PWL 0.1
`define FD4TQHSX4_CP_PWH 0.1
`define FD4TQHSX4_CP_PWL 0.1
`define FD4TQHSX4_D_CP_SETUP_posedge_posedge 0.1
`define FD4TQHSX4_D_CP_SETUP_negedge_posedge 0.1
`define FD4TQHSX4_D_CP_HOLD_posedge_posedge 0.1
`define FD4TQHSX4_D_CP_HOLD_negedge_posedge 0.1
`define FD4TQHSX4_TI_CP_SETUP_posedge_posedge 0.1
`define FD4TQHSX4_TI_CP_SETUP_negedge_posedge 0.1
`define FD4TQHSX4_TI_CP_HOLD_posedge_posedge 0.1
`define FD4TQHSX4_TI_CP_HOLD_negedge_posedge 0.1
`define FD4TQHSX4_TE_CP_SETUP_posedge_posedge 0.1
`define FD4TQHSX4_TE_CP_SETUP_negedge_posedge 0.1
`define FD4TQHSX4_TE_CP_HOLD_posedge_posedge 0.1
`define FD4TQHSX4_TE_CP_HOLD_negedge_posedge 0.1

module FD4TQHSX4 (Q, SO, D, CP, SD, TI, TE);

   output Q;
   output SO;
   input D;
   input CP;
   input SD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_FD_P_SN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, CP, SD, Notifier);

   buf  u2 (Q, IQ);
   buf  u3 (SO, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   and  (AndSDTEX_, SD, TEX);
   and  (AndSDTE_, SD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_SD_, XorDTI_, SD);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   nor  (D_orTI_onTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if(!TE && SD) (posedge CP => (Q +: D)) = (`FD4TQHSX4_CP_R_Q_R, `FD4TQHSX4_CP_R_Q_F);
      if(TE && SD) (posedge CP => (Q +: TI)) = (`FD4TQHSX4_CP_R_Q_R, `FD4TQHSX4_CP_R_Q_F);
      if(!D && TI && SD) (posedge CP => (Q +: TE)) = (`FD4TQHSX4_CP_R_Q_R, `FD4TQHSX4_CP_R_Q_F);
      if(!TI && D && SD) (posedge CP => (Q -: TE)) = (`FD4TQHSX4_CP_R_Q_R, `FD4TQHSX4_CP_R_Q_F);
      if(!TE && SD) (posedge CP => (SO +: D)) = (`FD4TQHSX4_CP_R_SO_R, `FD4TQHSX4_CP_R_SO_F);
      if(TE && SD) (posedge CP => (SO +: TI)) = (`FD4TQHSX4_CP_R_SO_R, `FD4TQHSX4_CP_R_SO_F);
      if(!D && TI && SD) (posedge CP => (SO +: TE)) = (`FD4TQHSX4_CP_R_SO_R, `FD4TQHSX4_CP_R_SO_F);
      if(!TI && D && SD) (posedge CP => (SO -: TE)) = (`FD4TQHSX4_CP_R_SO_R, `FD4TQHSX4_CP_R_SO_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4TQHSX4_SD_F_Q_R,`FD4TQHSX4_SD_F_Q_R);
      (negedge SD => (SO +: 1'b1)) = (`FD4TQHSX4_SD_F_SO_R,`FD4TQHSX4_SD_F_SO_R);

	$setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FD4TQHSX4_TE_CP_SETUP_posedge_posedge, `FD4TQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FD4TQHSX4_TE_CP_SETUP_negedge_posedge, `FD4TQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTE_, posedge TI, `FD4TQHSX4_TI_CP_SETUP_posedge_posedge, `FD4TQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTE_, negedge TI, `FD4TQHSX4_TI_CP_SETUP_negedge_posedge, `FD4TQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndSDTEX_, posedge D, `FD4TQHSX4_D_CP_SETUP_posedge_posedge, `FD4TQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndSDTEX_, negedge D, `FD4TQHSX4_D_CP_SETUP_negedge_posedge, `FD4TQHSX4_D_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD4TQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4TQHSX4_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4TQHSX4_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FD4TQHSX4_SD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& D_orTI_onTE, posedge SD, `FD4TQHSX4_SD_CP_REM_posedge_posedge, Notifier);
`else
       (posedge CP => (Q +: Mux21DTITE_)) = (`FD4TQHSX4_CP_R_Q_R, `FD4TQHSX4_CP_R_Q_F);
       (posedge CP => (SO +: Mux21DTITE_)) = (`FD4TQHSX4_CP_R_SO_R, `FD4TQHSX4_CP_R_SO_F);
      (negedge SD => (Q +: 1'b1)) = (`FD4TQHSX4_SD_F_Q_R,`FD4TQHSX4_SD_F_Q_R);
      (negedge SD => (SO +: 1'b1)) = (`FD4TQHSX4_SD_F_SO_R,`FD4TQHSX4_SD_F_SO_R);
 
        $setuphold(posedge CP &&& AndXorDTI_SD_, posedge TE, `FD4TQHSX4_TE_CP_SETUP_posedge_posedge, `FD4TQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndXorDTI_SD_, negedge TE, `FD4TQHSX4_TE_CP_SETUP_negedge_posedge, `FD4TQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTE_, posedge TI, `FD4TQHSX4_TI_CP_SETUP_posedge_posedge, `FD4TQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTE_, negedge TI, `FD4TQHSX4_TI_CP_SETUP_negedge_posedge, `FD4TQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndSDTEX_, posedge D, `FD4TQHSX4_D_CP_SETUP_posedge_posedge,`FD4TQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndSDTEX_, negedge D, `FD4TQHSX4_D_CP_SETUP_negedge_posedge,`FD4TQHSX4_D_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD4TQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP &&& SD, `FD4TQHSX4_CP_PWH, 0, Notifier);
      $width(negedge SD, `FD4TQHSX4_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& D_orTI_onTE, `FD4TQHSX4_SD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& D_orTI_onTE, posedge SD, `FD4TQHSX4_SD_CP_REM_posedge_posedge, Notifier);

`endif

   endspecify
`endif


endmodule // FD4TQHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:44 and Version :1.1 //
 
//  START 
// CELL FD6SHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD6SHS_CP_R_QN_F 0.1
`define FD6SHS_CP_R_QN_R 0.1
`define FD6SHS_CP_R_Q_R 0.1
`define FD6SHS_CP_R_Q_F 0.1
`define FD6SHS_CP_PWH 0.1
`define FD6SHS_CP_PWL 0.1
`define FD6SHS_TE_CP_SETUP_posedge_posedge 0.1
`define FD6SHS_TE_CP_SETUP_negedge_posedge 0.1
`define FD6SHS_TE_CP_HOLD_posedge_posedge 0.1
`define FD6SHS_TE_CP_HOLD_negedge_posedge 0.1
`define FD6SHS_TI_CP_SETUP_posedge_posedge 0.1
`define FD6SHS_TI_CP_SETUP_negedge_posedge 0.1
`define FD6SHS_TI_CP_HOLD_posedge_posedge 0.1
`define FD6SHS_TI_CP_HOLD_negedge_posedge 0.1
`define FD6SHS_S_CP_SETUP_posedge_posedge 0.1
`define FD6SHS_S_CP_SETUP_negedge_posedge 0.1
`define FD6SHS_S_CP_HOLD_posedge_posedge 0.1
`define FD6SHS_S_CP_HOLD_negedge_posedge 0.1
`define FD6SHS_D0_CP_SETUP_posedge_posedge 0.1
`define FD6SHS_D0_CP_SETUP_negedge_posedge 0.1
`define FD6SHS_D0_CP_HOLD_posedge_posedge 0.1
`define FD6SHS_D0_CP_HOLD_negedge_posedge 0.1
`define FD6SHS_D1_CP_SETUP_posedge_posedge 0.1
`define FD6SHS_D1_CP_SETUP_negedge_posedge 0.1
`define FD6SHS_D1_CP_HOLD_posedge_posedge 0.1
`define FD6SHS_D1_CP_HOLD_negedge_posedge 0.1

module FD6SHS (Q, QN, D0, D1, S, CP, TI, TE);

   output Q;
   output QN;
   input CP;
   input TE;
   input TI;
   input S;
   input D0;
   input D1;


   reg Notifier;

   U_MUX2  u0 (Mux21D0D1S_, D0, D1, S);
   U_MUX2  u1 (Mux21Mux21D0D1S_TITE_, Mux21D0D1S_, TI, TE);

   U_FD_P_NOTI u2 (   // Verilog Seq UDP
      IQ, Mux21Mux21D0D1S_TITE_, CP, Notifier);

   buf  u3 (Q, IQ);
   not  u4 (QN, IQ);



`ifdef functional
`else
   xor  (D_orTI, Mux21D0D1S_, TI);
   not  (SX, S);
   not  (TIX, TI);
   not  (D1X, D1);
   or  (OrTED0D1X_, TE, D0, D1X);
   not  (D0X, D0);
   or  (OrTED0XD1_, TE, D0X, D1);
   nand  (NandOrTED0D1X_OrTED0XD1__, OrTED0D1X_, OrTED0XD1_);
   nor  (NorTES_, TE, S);
   not  (TEX, TE);
   and  (AndTEXS_, TEX, S);
   specify
`ifdef verifault

      if(!D0 && !S && TI) (posedge CP => (Q +: TE)) = (`FD6SHS_CP_R_Q_R, `FD6SHS_CP_R_Q_F);
      if(!D1 && S && TI) (posedge CP => (Q +: TE)) = (`FD6SHS_CP_R_Q_R, `FD6SHS_CP_R_Q_F);
      if(!TI && S && D1) (posedge CP => (Q -: TE)) = (`FD6SHS_CP_R_Q_R, `FD6SHS_CP_R_Q_F);
      if(!TI && !S && D0) (posedge CP => (Q -: TE)) = (`FD6SHS_CP_R_Q_R, `FD6SHS_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD6SHS_CP_R_Q_R, `FD6SHS_CP_R_Q_F);
      if(!D0 && !TE && D1) (posedge CP => (Q +: S)) = (`FD6SHS_CP_R_Q_R, `FD6SHS_CP_R_Q_F);
      if(!D1 && !TE && D0) (posedge CP => (Q -: S)) = (`FD6SHS_CP_R_Q_R, `FD6SHS_CP_R_Q_F);
      if(!TE && !S) (posedge CP => (Q +: D0)) = (`FD6SHS_CP_R_Q_R, `FD6SHS_CP_R_Q_F);
      if(!TE && S) (posedge CP => (Q +: D1)) = (`FD6SHS_CP_R_Q_R, `FD6SHS_CP_R_Q_F);
      if(!D0 && !S && TI) (posedge CP => (QN -: TE)) = (`FD6SHS_CP_R_QN_R, `FD6SHS_CP_R_QN_F);
      if(!D1 && S && TI) (posedge CP => (QN -: TE)) = (`FD6SHS_CP_R_QN_R, `FD6SHS_CP_R_QN_F);
      if(!TI && S && D1) (posedge CP => (QN +: TE)) = (`FD6SHS_CP_R_QN_R, `FD6SHS_CP_R_QN_F);
      if(!TI && !S && D0) (posedge CP => (QN +: TE)) = (`FD6SHS_CP_R_QN_R, `FD6SHS_CP_R_QN_F);
      if(TE) (posedge CP => (QN -: TI)) = (`FD6SHS_CP_R_QN_R, `FD6SHS_CP_R_QN_F);
      if(!D0 && !TE && D1) (posedge CP => (QN -: S)) = (`FD6SHS_CP_R_QN_R, `FD6SHS_CP_R_QN_F);
      if(!D1 && !TE && D0) (posedge CP => (QN +: S)) = (`FD6SHS_CP_R_QN_R, `FD6SHS_CP_R_QN_F);
      if(!TE && !S) (posedge CP => (QN -: D0)) = (`FD6SHS_CP_R_QN_R, `FD6SHS_CP_R_QN_F);
      if(!TE && S) (posedge CP => (QN -: D1)) = (`FD6SHS_CP_R_QN_R, `FD6SHS_CP_R_QN_F);

	$setuphold(posedge CP &&& AndTEXS_, posedge D1, `FD6SHS_D1_CP_SETUP_posedge_posedge, `FD6SHS_D1_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndTEXS_, negedge D1, `FD6SHS_D1_CP_SETUP_negedge_posedge, `FD6SHS_D1_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& NorTES_, posedge D0, `FD6SHS_D0_CP_SETUP_posedge_posedge, `FD6SHS_D0_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& NorTES_, negedge D0, `FD6SHS_D0_CP_SETUP_negedge_posedge, `FD6SHS_D0_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& NandOrTED0D1X_OrTED0XD1__, posedge S, `FD6SHS_S_CP_SETUP_posedge_posedge, `FD6SHS_S_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& NandOrTED0D1X_OrTED0XD1__, negedge S, `FD6SHS_S_CP_SETUP_negedge_posedge, `FD6SHS_S_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FD6SHS_TI_CP_SETUP_posedge_posedge, `FD6SHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FD6SHS_TI_CP_SETUP_negedge_posedge, `FD6SHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& D_orTI, posedge TE, `FD6SHS_TE_CP_SETUP_posedge_posedge, `FD6SHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& D_orTI, negedge TE, `FD6SHS_TE_CP_SETUP_negedge_posedge, `FD6SHS_TE_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD6SHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD6SHS_CP_PWH, 0, Notifier);
`else
      (posedge CP => (Q +: Mux21Mux21D0D1S_TITE_)) = (`FD6SHS_CP_R_Q_R, `FD6SHS_CP_R_Q_F);
      (posedge CP => (QN -: Mux21Mux21D0D1S_TITE_)) = (`FD6SHS_CP_R_QN_R, `FD6SHS_CP_R_QN_F);
 
        $setuphold(posedge CP &&& AndTEXS_, posedge D1, `FD6SHS_D1_CP_SETUP_posedge_posedge,`FD6SHS_D1_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndTEXS_, negedge D1, `FD6SHS_D1_CP_SETUP_negedge_posedge,`FD6SHS_D1_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& NorTES_, posedge D0, `FD6SHS_D0_CP_SETUP_posedge_posedge,`FD6SHS_D0_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& NorTES_, negedge D0, `FD6SHS_D0_CP_SETUP_negedge_posedge,`FD6SHS_D0_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& NandOrTED0D1X_OrTED0XD1__, posedge S, `FD6SHS_S_CP_SETUP_posedge_posedge, `FD6SHS_S_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& NandOrTED0D1X_OrTED0XD1__, negedge S, `FD6SHS_S_CP_SETUP_negedge_posedge, `FD6SHS_S_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD6SHS_TI_CP_SETUP_posedge_posedge, `FD6SHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD6SHS_TI_CP_SETUP_negedge_posedge, `FD6SHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& D_orTI, posedge TE, `FD6SHS_TE_CP_SETUP_posedge_posedge, `FD6SHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& D_orTI, negedge TE, `FD6SHS_TE_CP_SETUP_negedge_posedge, `FD6SHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD6SHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD6SHS_CP_PWH, 0, Notifier);
`endif
   endspecify
`endif


endmodule // FD6SHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:50 and Version :1.1 //
 
//  START 
// CELL FD6SQHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD6SQHS_CP_R_Q_R 0.1
`define FD6SQHS_CP_R_Q_F 0.1
`define FD6SQHS_CP_PWH 0.1
`define FD6SQHS_CP_PWL 0.1
`define FD6SQHS_TE_CP_SETUP_posedge_posedge 0.1
`define FD6SQHS_TE_CP_SETUP_negedge_posedge 0.1
`define FD6SQHS_TE_CP_HOLD_posedge_posedge 0.1
`define FD6SQHS_TE_CP_HOLD_negedge_posedge 0.1
`define FD6SQHS_TI_CP_SETUP_posedge_posedge 0.1
`define FD6SQHS_TI_CP_SETUP_negedge_posedge 0.1
`define FD6SQHS_TI_CP_HOLD_posedge_posedge 0.1
`define FD6SQHS_TI_CP_HOLD_negedge_posedge 0.1
`define FD6SQHS_S_CP_SETUP_posedge_posedge 0.1
`define FD6SQHS_S_CP_SETUP_negedge_posedge 0.1
`define FD6SQHS_S_CP_HOLD_posedge_posedge 0.1
`define FD6SQHS_S_CP_HOLD_negedge_posedge 0.1
`define FD6SQHS_D0_CP_SETUP_posedge_posedge 0.1
`define FD6SQHS_D0_CP_SETUP_negedge_posedge 0.1
`define FD6SQHS_D0_CP_HOLD_posedge_posedge 0.1
`define FD6SQHS_D0_CP_HOLD_negedge_posedge 0.1
`define FD6SQHS_D1_CP_SETUP_posedge_posedge 0.1
`define FD6SQHS_D1_CP_SETUP_negedge_posedge 0.1
`define FD6SQHS_D1_CP_HOLD_posedge_posedge 0.1
`define FD6SQHS_D1_CP_HOLD_negedge_posedge 0.1

module FD6SQHS (Q, D0, D1, S, CP, TI, TE);

   output Q;
   input CP;
   input TE;
   input TI;
   input S;
   input D0;
   input D1;


   reg Notifier;

   U_MUX2  u0 (Mux21D0D1S_, D0, D1, S);
   U_MUX2  u1 (Mux21Mux21D0D1S_TITE_, Mux21D0D1S_, TI, TE);

   U_FD_P_NOTI u2 (   // Verilog Seq UDP
      IQ, Mux21Mux21D0D1S_TITE_, CP, Notifier);

   buf  u3 (Q, IQ);



`ifdef functional
`else
   xor  (D_orTI, Mux21D0D1S_, TI);
   not  (SX, S);
   not  (TIX, TI);
   not  (D1X, D1);
   or  (OrTED0D1X_, TE, D0, D1X);
   not  (D0X, D0);
   or  (OrTED0XD1_, TE, D0X, D1);
   nand  (NandOrTED0D1X_OrTED0XD1__, OrTED0D1X_, OrTED0XD1_);
   nor  (NorTES_, TE, S);
   not  (TEX, TE);
   and  (AndTEXS_, TEX, S);
   specify
`ifdef verifault 

      if(!D0 && !S && TI) (posedge CP => (Q +: TE)) = (`FD6SQHS_CP_R_Q_R, `FD6SQHS_CP_R_Q_F);
      if(!D1 && S && TI) (posedge CP => (Q +: TE)) = (`FD6SQHS_CP_R_Q_R, `FD6SQHS_CP_R_Q_F);
      if(!TI && S && D1) (posedge CP => (Q -: TE)) = (`FD6SQHS_CP_R_Q_R, `FD6SQHS_CP_R_Q_F);
      if(!TI && !S && D0) (posedge CP => (Q -: TE)) = (`FD6SQHS_CP_R_Q_R, `FD6SQHS_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD6SQHS_CP_R_Q_R, `FD6SQHS_CP_R_Q_F);
      if(!D0 && !TE && D1) (posedge CP => (Q +: S)) = (`FD6SQHS_CP_R_Q_R, `FD6SQHS_CP_R_Q_F);
      if(!D1 && !TE && D0) (posedge CP => (Q -: S)) = (`FD6SQHS_CP_R_Q_R, `FD6SQHS_CP_R_Q_F);
      if(!TE && !S) (posedge CP => (Q +: D0)) = (`FD6SQHS_CP_R_Q_R, `FD6SQHS_CP_R_Q_F);
      if(!TE && S) (posedge CP => (Q +: D1)) = (`FD6SQHS_CP_R_Q_R, `FD6SQHS_CP_R_Q_F);

	$setuphold(posedge CP &&& AndTEXS_, posedge D1, `FD6SQHS_D1_CP_SETUP_posedge_posedge, `FD6SQHS_D1_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndTEXS_, negedge D1, `FD6SQHS_D1_CP_SETUP_negedge_posedge, `FD6SQHS_D1_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& NorTES_, posedge D0, `FD6SQHS_D0_CP_SETUP_posedge_posedge, `FD6SQHS_D0_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& NorTES_, negedge D0, `FD6SQHS_D0_CP_SETUP_negedge_posedge, `FD6SQHS_D0_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& NandOrTED0D1X_OrTED0XD1__, posedge S, `FD6SQHS_S_CP_SETUP_posedge_posedge, `FD6SQHS_S_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& NandOrTED0D1X_OrTED0XD1__, negedge S, `FD6SQHS_S_CP_SETUP_negedge_posedge, `FD6SQHS_S_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FD6SQHS_TI_CP_SETUP_posedge_posedge, `FD6SQHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FD6SQHS_TI_CP_SETUP_negedge_posedge, `FD6SQHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& D_orTI, posedge TE, `FD6SQHS_TE_CP_SETUP_posedge_posedge, `FD6SQHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& D_orTI, negedge TE, `FD6SQHS_TE_CP_SETUP_negedge_posedge, `FD6SQHS_TE_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD6SQHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD6SQHS_CP_PWH, 0, Notifier);
`else
      (posedge CP => (Q +: Mux21Mux21D0D1S_TITE_)) = (`FD6SQHS_CP_R_Q_R, `FD6SQHS_CP_R_Q_F);
 
        $setuphold(posedge CP &&& AndTEXS_, posedge D1, `FD6SQHS_D1_CP_SETUP_posedge_posedge, `FD6SQHS_D1_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndTEXS_, negedge D1, `FD6SQHS_D1_CP_SETUP_negedge_posedge, `FD6SQHS_D1_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& NorTES_, posedge D0, `FD6SQHS_D0_CP_SETUP_posedge_posedge, `FD6SQHS_D0_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& NorTES_, negedge D0, `FD6SQHS_D0_CP_SETUP_negedge_posedge, `FD6SQHS_D0_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& NandOrTED0D1X_OrTED0XD1__, posedge S, `FD6SQHS_S_CP_SETUP_posedge_posedge, `FD6SQHS_S_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& NandOrTED0D1X_OrTED0XD1__, negedge S, `FD6SQHS_S_CP_SETUP_negedge_posedge, `FD6SQHS_S_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD6SQHS_TI_CP_SETUP_posedge_posedge, `FD6SQHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD6SQHS_TI_CP_SETUP_negedge_posedge, `FD6SQHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& D_orTI, posedge TE, `FD6SQHS_TE_CP_SETUP_posedge_posedge, `FD6SQHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& D_orTI, negedge TE, `FD6SQHS_TE_CP_SETUP_negedge_posedge, `FD6SQHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD6SQHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD6SQHS_CP_PWH, 0, Notifier);
`endif

   endspecify
`endif


endmodule // FD6SQHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:54 and Version :1.1 //
 
//  START 
// CELL FD6THS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD6THS_CP_R_QN_F 0.1
`define FD6THS_CP_R_QN_R 0.1
`define FD6THS_CP_R_Q_R 0.1
`define FD6THS_CP_R_Q_F 0.1
`define FD6THS_CP_R_SO_R 0.1
`define FD6THS_CP_R_SO_F 0.1
`define FD6THS_CP_PWH 0.1
`define FD6THS_CP_PWL 0.1
`define FD6THS_TE_CP_SETUP_posedge_posedge 0.1
`define FD6THS_TE_CP_SETUP_negedge_posedge 0.1
`define FD6THS_TE_CP_HOLD_posedge_posedge 0.1
`define FD6THS_TE_CP_HOLD_negedge_posedge 0.1
`define FD6THS_TI_CP_SETUP_posedge_posedge 0.1
`define FD6THS_TI_CP_SETUP_negedge_posedge 0.1
`define FD6THS_TI_CP_HOLD_posedge_posedge 0.1
`define FD6THS_TI_CP_HOLD_negedge_posedge 0.1
`define FD6THS_S_CP_SETUP_posedge_posedge 0.1
`define FD6THS_S_CP_SETUP_negedge_posedge 0.1
`define FD6THS_S_CP_HOLD_posedge_posedge 0.1
`define FD6THS_S_CP_HOLD_negedge_posedge 0.1
`define FD6THS_D0_CP_SETUP_posedge_posedge 0.1
`define FD6THS_D0_CP_SETUP_negedge_posedge 0.1
`define FD6THS_D0_CP_HOLD_posedge_posedge 0.1
`define FD6THS_D0_CP_HOLD_negedge_posedge 0.1
`define FD6THS_D1_CP_SETUP_posedge_posedge 0.1
`define FD6THS_D1_CP_SETUP_negedge_posedge 0.1
`define FD6THS_D1_CP_HOLD_posedge_posedge 0.1
`define FD6THS_D1_CP_HOLD_negedge_posedge 0.1

module FD6THS (Q, QN, SO, D0, D1, S, CP, TI, TE);

   output Q;
   output QN;
   output SO;
   input CP;
   input TE;
   input TI;
   input S;
   input D0;
   input D1;


   reg Notifier;

   U_MUX2  u0 (Mux21D0D1S_, D0, D1, S);
   U_MUX2  u1 (Mux21Mux21D0D1S_TITE_, Mux21D0D1S_, TI, TE);

   U_FD_P_NOTI u2 (   // Verilog Seq UDP
      IQ, Mux21Mux21D0D1S_TITE_, CP, Notifier);

   buf  u3 (Q, IQ);
   not  u4 (QN, IQ);
   buf  u5 (SO, IQ);



`ifdef functional
`else
   xor  (D_orTI, Mux21D0D1S_, TI);
   not  (SX, S);
   not  (TIX, TI);
   not  (D1X, D1);
   or  (OrTED0D1X_, TE, D0, D1X);
   not  (D0X, D0);
   or  (OrTED0XD1_, TE, D0X, D1);
   nand  (NandOrTED0D1X_OrTED0XD1__, OrTED0D1X_, OrTED0XD1_);
   nor  (NorTES_, TE, S);
   not  (TEX, TE);
   and  (AndTEXS_, TEX, S);
   specify
`ifdef verifault

      if(!D0 && !S && TI) (posedge CP => (Q +: TE)) = (`FD6THS_CP_R_Q_R, `FD6THS_CP_R_Q_F);
      if(!D1 && S && TI) (posedge CP => (Q +: TE)) = (`FD6THS_CP_R_Q_R, `FD6THS_CP_R_Q_F);
      if(!TI && S && D1) (posedge CP => (Q -: TE)) = (`FD6THS_CP_R_Q_R, `FD6THS_CP_R_Q_F);
      if(!TI && !S && D0) (posedge CP => (Q -: TE)) = (`FD6THS_CP_R_Q_R, `FD6THS_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD6THS_CP_R_Q_R, `FD6THS_CP_R_Q_F);
      if(!D0 && !TE && D1) (posedge CP => (Q +: S)) = (`FD6THS_CP_R_Q_R, `FD6THS_CP_R_Q_F);
      if(!D1 && !TE && D0) (posedge CP => (Q -: S)) = (`FD6THS_CP_R_Q_R, `FD6THS_CP_R_Q_F);
      if(!TE && !S) (posedge CP => (Q +: D0)) = (`FD6THS_CP_R_Q_R, `FD6THS_CP_R_Q_F);
      if(!TE && S) (posedge CP => (Q +: D1)) = (`FD6THS_CP_R_Q_R, `FD6THS_CP_R_Q_F);
      if(!D0 && !S && TI) (posedge CP => (QN -: TE)) = (`FD6THS_CP_R_QN_R, `FD6THS_CP_R_QN_F);
      if(!D1 && S && TI) (posedge CP => (QN -: TE)) = (`FD6THS_CP_R_QN_R, `FD6THS_CP_R_QN_F);
      if(!TI && S && D1) (posedge CP => (QN +: TE)) = (`FD6THS_CP_R_QN_R, `FD6THS_CP_R_QN_F);
      if(!TI && !S && D0) (posedge CP => (QN +: TE)) = (`FD6THS_CP_R_QN_R, `FD6THS_CP_R_QN_F);
      if(TE) (posedge CP => (QN -: TI)) = (`FD6THS_CP_R_QN_R, `FD6THS_CP_R_QN_F);
      if(!D0 && !TE && D1) (posedge CP => (QN -: S)) = (`FD6THS_CP_R_QN_R, `FD6THS_CP_R_QN_F);
      if(!D1 && !TE && D0) (posedge CP => (QN +: S)) = (`FD6THS_CP_R_QN_R, `FD6THS_CP_R_QN_F);
      if(!TE && !S) (posedge CP => (QN -: D0)) = (`FD6THS_CP_R_QN_R, `FD6THS_CP_R_QN_F);
      if(!TE && S) (posedge CP => (QN -: D1)) = (`FD6THS_CP_R_QN_R, `FD6THS_CP_R_QN_F);

      if(!D0 && !S && TI) (posedge CP => (SO +: TE)) = (`FD6THS_CP_R_SO_R, `FD6THS_CP_R_SO_F);
      if(!D1 && S && TI) (posedge CP => (SO +: TE)) = (`FD6THS_CP_R_SO_R, `FD6THS_CP_R_SO_F);
      if(!TI && S && D1) (posedge CP => (SO -: TE)) = (`FD6THS_CP_R_SO_R, `FD6THS_CP_R_SO_F);
      if(!TI && !S && D0) (posedge CP => (SO -: TE)) = (`FD6THS_CP_R_SO_R, `FD6THS_CP_R_SO_F);
      if(TE) (posedge CP => (SO +: TI)) = (`FD6THS_CP_R_SO_R, `FD6THS_CP_R_SO_F);
      if(!D0 && !TE && D1) (posedge CP => (SO +: S)) = (`FD6THS_CP_R_SO_R, `FD6THS_CP_R_SO_F);
      if(!D1 && !TE && D0) (posedge CP => (SO -: S)) = (`FD6THS_CP_R_SO_R, `FD6THS_CP_R_SO_F);
      if(!TE && !S) (posedge CP => (SO +: D0)) = (`FD6THS_CP_R_SO_R, `FD6THS_CP_R_SO_F);
      if(!TE && S) (posedge CP => (SO +: D1)) = (`FD6THS_CP_R_SO_R, `FD6THS_CP_R_SO_F);

	$setuphold(posedge CP &&& AndTEXS_, posedge D1, `FD6THS_D1_CP_SETUP_posedge_posedge, `FD6THS_D1_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndTEXS_, negedge D1, `FD6THS_D1_CP_SETUP_negedge_posedge, `FD6THS_D1_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& NorTES_, posedge D0, `FD6THS_D0_CP_SETUP_posedge_posedge, `FD6THS_D0_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& NorTES_, negedge D0, `FD6THS_D0_CP_SETUP_negedge_posedge, `FD6THS_D0_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& NandOrTED0D1X_OrTED0XD1__, posedge S, `FD6THS_S_CP_SETUP_posedge_posedge, `FD6THS_S_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& NandOrTED0D1X_OrTED0XD1__, negedge S, `FD6THS_S_CP_SETUP_negedge_posedge, `FD6THS_S_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FD6THS_TI_CP_SETUP_posedge_posedge, `FD6THS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FD6THS_TI_CP_SETUP_negedge_posedge, `FD6THS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& D_orTI, posedge TE, `FD6THS_TE_CP_SETUP_posedge_posedge, `FD6THS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& D_orTI, negedge TE, `FD6THS_TE_CP_SETUP_negedge_posedge, `FD6THS_TE_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD6THS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD6THS_CP_PWH, 0, Notifier);
`else

      (posedge CP => (Q +: Mux21Mux21D0D1S_TITE_)) = (`FD6THS_CP_R_Q_R, `FD6THS_CP_R_Q_F);
      (posedge CP => (QN -: Mux21Mux21D0D1S_TITE_)) = (`FD6THS_CP_R_QN_R, `FD6THS_CP_R_QN_F);
 
      (posedge CP => (SO +: Mux21Mux21D0D1S_TITE_)) = (`FD6THS_CP_R_SO_R, `FD6THS_CP_R_SO_F);
 
        $setuphold(posedge CP &&& AndTEXS_, posedge D1, `FD6THS_D1_CP_SETUP_posedge_posedge, `FD6THS_D1_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndTEXS_, negedge D1, `FD6THS_D1_CP_SETUP_negedge_posedge, `FD6THS_D1_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& NorTES_, posedge D0, `FD6THS_D0_CP_SETUP_posedge_posedge, `FD6THS_D0_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& NorTES_, negedge D0, `FD6THS_D0_CP_SETUP_negedge_posedge, `FD6THS_D0_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& NandOrTED0D1X_OrTED0XD1__, posedge S, `FD6THS_S_CP_SETUP_posedge_posedge, `FD6THS_S_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& NandOrTED0D1X_OrTED0XD1__, negedge S, `FD6THS_S_CP_SETUP_negedge_posedge, `FD6THS_S_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD6THS_TI_CP_SETUP_posedge_posedge, `FD6THS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD6THS_TI_CP_SETUP_negedge_posedge, `FD6THS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& D_orTI, posedge TE, `FD6THS_TE_CP_SETUP_posedge_posedge, `FD6THS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& D_orTI, negedge TE, `FD6THS_TE_CP_SETUP_negedge_posedge, `FD6THS_TE_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD6THS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD6THS_CP_PWH, 0, Notifier);
`endif
   endspecify
`endif


endmodule // FD6THS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:50 and Version :1.1 //
 
//  START 
// CELL FD6TQHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD6TQHS_CP_R_Q_R 0.1
`define FD6TQHS_CP_R_Q_F 0.1
`define FD6TQHS_CP_R_SO_R 0.1
`define FD6TQHS_CP_R_SO_F 0.1
`define FD6TQHS_CP_PWH 0.1
`define FD6TQHS_CP_PWL 0.1
`define FD6TQHS_TE_CP_SETUP_posedge_posedge 0.1
`define FD6TQHS_TE_CP_SETUP_negedge_posedge 0.1
`define FD6TQHS_TE_CP_HOLD_posedge_posedge 0.1
`define FD6TQHS_TE_CP_HOLD_negedge_posedge 0.1
`define FD6TQHS_TI_CP_SETUP_posedge_posedge 0.1
`define FD6TQHS_TI_CP_SETUP_negedge_posedge 0.1
`define FD6TQHS_TI_CP_HOLD_posedge_posedge 0.1
`define FD6TQHS_TI_CP_HOLD_negedge_posedge 0.1
`define FD6TQHS_S_CP_SETUP_posedge_posedge 0.1
`define FD6TQHS_S_CP_SETUP_negedge_posedge 0.1
`define FD6TQHS_S_CP_HOLD_posedge_posedge 0.1
`define FD6TQHS_S_CP_HOLD_negedge_posedge 0.1
`define FD6TQHS_D0_CP_SETUP_posedge_posedge 0.1
`define FD6TQHS_D0_CP_SETUP_negedge_posedge 0.1
`define FD6TQHS_D0_CP_HOLD_posedge_posedge 0.1
`define FD6TQHS_D0_CP_HOLD_negedge_posedge 0.1
`define FD6TQHS_D1_CP_SETUP_posedge_posedge 0.1
`define FD6TQHS_D1_CP_SETUP_negedge_posedge 0.1
`define FD6TQHS_D1_CP_HOLD_posedge_posedge 0.1
`define FD6TQHS_D1_CP_HOLD_negedge_posedge 0.1

module FD6TQHS (Q, SO, D0, D1, S, CP, TI, TE);

   output Q;
   output SO;
   input CP;
   input TE;
   input TI;
   input S;
   input D0;
   input D1;


   reg Notifier;

   U_MUX2  u0 (Mux21D0D1S_, D0, D1, S);
   U_MUX2  u1 (Mux21Mux21D0D1S_TITE_, Mux21D0D1S_, TI, TE);

   U_FD_P_NOTI u2 (   // Verilog Seq UDP
      IQ, Mux21Mux21D0D1S_TITE_, CP, Notifier);

   buf  u3 (Q, IQ);
   buf  u5 (SO, IQ);



`ifdef functional
`else
   xor  (D_orTI, Mux21D0D1S_, TI);
   not  (SX, S);
   not  (TIX, TI);
   not  (D1X, D1);
   or  (OrTED0D1X_, TE, D0, D1X);
   not  (D0X, D0);
   or  (OrTED0XD1_, TE, D0X, D1);
   nand  (NandOrTED0D1X_OrTED0XD1__, OrTED0D1X_, OrTED0XD1_);
   nor  (NorTES_, TE, S);
   not  (TEX, TE);
   and  (AndTEXS_, TEX, S);
   specify
`ifdef verifault

      if(!D0 && !S && TI) (posedge CP => (Q +: TE)) = (`FD6TQHS_CP_R_Q_R, `FD6TQHS_CP_R_Q_F);
      if(!D1 && S && TI) (posedge CP => (Q +: TE)) = (`FD6TQHS_CP_R_Q_R, `FD6TQHS_CP_R_Q_F);
      if(!TI && S && D1) (posedge CP => (Q -: TE)) = (`FD6TQHS_CP_R_Q_R, `FD6TQHS_CP_R_Q_F);
      if(!TI && !S && D0) (posedge CP => (Q -: TE)) = (`FD6TQHS_CP_R_Q_R, `FD6TQHS_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD6TQHS_CP_R_Q_R, `FD6TQHS_CP_R_Q_F);
      if(!D0 && !TE && D1) (posedge CP => (Q +: S)) = (`FD6TQHS_CP_R_Q_R, `FD6TQHS_CP_R_Q_F);
      if(!D1 && !TE && D0) (posedge CP => (Q -: S)) = (`FD6TQHS_CP_R_Q_R, `FD6TQHS_CP_R_Q_F);
      if(!TE && !S) (posedge CP => (Q +: D0)) = (`FD6TQHS_CP_R_Q_R, `FD6TQHS_CP_R_Q_F);
      if(!TE && S) (posedge CP => (Q +: D1)) = (`FD6TQHS_CP_R_Q_R, `FD6TQHS_CP_R_Q_F);

      if(!D0 && !S && TI) (posedge CP => (SO +: TE)) = (`FD6TQHS_CP_R_SO_R, `FD6TQHS_CP_R_SO_F);
      if(!D1 && S && TI) (posedge CP => (SO +: TE)) = (`FD6TQHS_CP_R_SO_R, `FD6TQHS_CP_R_SO_F);
      if(!TI && S && D1) (posedge CP => (SO -: TE)) = (`FD6TQHS_CP_R_SO_R, `FD6TQHS_CP_R_SO_F);
      if(!TI && !S && D0) (posedge CP => (SO -: TE)) = (`FD6TQHS_CP_R_SO_R, `FD6TQHS_CP_R_SO_F);
      if(TE) (posedge CP => (SO +: TI)) = (`FD6TQHS_CP_R_SO_R, `FD6TQHS_CP_R_SO_F);
      if(!D0 && !TE && D1) (posedge CP => (SO +: S)) = (`FD6TQHS_CP_R_SO_R, `FD6TQHS_CP_R_SO_F);
      if(!D1 && !TE && D0) (posedge CP => (SO -: S)) = (`FD6TQHS_CP_R_SO_R, `FD6TQHS_CP_R_SO_F);
      if(!TE && !S) (posedge CP => (SO +: D0)) = (`FD6TQHS_CP_R_SO_R, `FD6TQHS_CP_R_SO_F);
      if(!TE && S) (posedge CP => (SO +: D1)) = (`FD6TQHS_CP_R_SO_R, `FD6TQHS_CP_R_SO_F);

	$setuphold(posedge CP &&& AndTEXS_, posedge D1, `FD6TQHS_D1_CP_SETUP_posedge_posedge, `FD6TQHS_D1_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndTEXS_, negedge D1, `FD6TQHS_D1_CP_SETUP_negedge_posedge, `FD6TQHS_D1_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& NorTES_, posedge D0, `FD6TQHS_D0_CP_SETUP_posedge_posedge, `FD6TQHS_D0_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& NorTES_, negedge D0, `FD6TQHS_D0_CP_SETUP_negedge_posedge, `FD6TQHS_D0_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& NandOrTED0D1X_OrTED0XD1__, posedge S, `FD6TQHS_S_CP_SETUP_posedge_posedge, `FD6TQHS_S_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& NandOrTED0D1X_OrTED0XD1__, negedge S, `FD6TQHS_S_CP_SETUP_negedge_posedge, `FD6TQHS_S_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FD6TQHS_TI_CP_SETUP_posedge_posedge, `FD6TQHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FD6TQHS_TI_CP_SETUP_negedge_posedge, `FD6TQHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& D_orTI, posedge TE, `FD6TQHS_TE_CP_SETUP_posedge_posedge, `FD6TQHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& D_orTI, negedge TE, `FD6TQHS_TE_CP_SETUP_negedge_posedge, `FD6TQHS_TE_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD6TQHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD6TQHS_CP_PWH, 0, Notifier);
`else
      (posedge CP => (Q +: Mux21Mux21D0D1S_TITE_)) = (`FD6TQHS_CP_R_Q_R, `FD6TQHS_CP_R_Q_F);
 
      (posedge CP => (SO +: Mux21Mux21D0D1S_TITE_)) = (`FD6TQHS_CP_R_SO_R, `FD6TQHS_CP_R_SO_F);
 
        $setuphold(posedge CP &&& AndTEXS_, posedge D1, `FD6TQHS_D1_CP_SETUP_posedge_posedge, `FD6TQHS_D1_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndTEXS_, negedge D1, `FD6TQHS_D1_CP_SETUP_negedge_posedge, `FD6TQHS_D1_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& NorTES_, posedge D0, `FD6TQHS_D0_CP_SETUP_posedge_posedge, `FD6TQHS_D0_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& NorTES_, negedge D0, `FD6TQHS_D0_CP_SETUP_negedge_posedge, `FD6TQHS_D0_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& NandOrTED0D1X_OrTED0XD1__, posedge S, `FD6TQHS_S_CP_SETUP_posedge_posedge, `FD6TQHS_S_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& NandOrTED0D1X_OrTED0XD1__, negedge S, `FD6TQHS_S_CP_SETUP_negedge_posedge, `FD6TQHS_S_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD6TQHS_TI_CP_SETUP_posedge_posedge, `FD6TQHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD6TQHS_TI_CP_SETUP_negedge_posedge, `FD6TQHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& D_orTI, posedge TE, `FD6TQHS_TE_CP_SETUP_posedge_posedge, `FD6TQHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& D_orTI, negedge TE, `FD6TQHS_TE_CP_SETUP_negedge_posedge, `FD6TQHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD6TQHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD6TQHS_CP_PWH, 0, Notifier);
 
`endif
   endspecify
`endif


endmodule // FD6TQHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:54 and Version :1.1 //
 
//  START 
// CELL FD7HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD7HS_CP_R_QN_F 0.1
`define FD7HS_CP_R_QN_R 0.1
`define FD7HS_CP_R_Q_R 0.1
`define FD7HS_CP_R_Q_F 0.1
`define FD7HS_CP_PWH 0.1
`define FD7HS_CP_PWL 0.1
`define FD7HS_E_CP_SETUP_posedge_posedge 0.1
`define FD7HS_E_CP_SETUP_negedge_posedge 0.1
`define FD7HS_E_CP_HOLD_posedge_posedge 0.1
`define FD7HS_E_CP_HOLD_negedge_posedge 0.1
`define FD7HS_D_CP_SETUP_posedge_posedge 0.1
`define FD7HS_D_CP_SETUP_negedge_posedge 0.1
`define FD7HS_D_CP_HOLD_posedge_posedge 0.1
`define FD7HS_D_CP_HOLD_negedge_posedge 0.1
 
module FD7HS (Q, QN, D, E, CP);
 
   output Q;
   output QN;
   input D;
   input E;
   input CP;
 
 
   reg Notifier;
 
   U_MUX2  u0 (Mux21IQDE_, IQ, D, E);
 
   U_FD_P_NOTI u2 (   // Verilog Seq UDP
     IQ, Mux21IQDE_, CP, Notifier);
 
   buf  u3 (Q, IQ);
   not  u4 (QN, IQ);
 
 
 
`ifdef functional
`else
   specify
 
      (posedge CP => (Q +: D)) = (`FD7HS_CP_R_Q_R, `FD7HS_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`FD7HS_CP_R_QN_R, `FD7HS_CP_R_QN_F);
 
	$setuphold(posedge CP &&& E, posedge D, `FD7HS_D_CP_SETUP_posedge_posedge, `FD7HS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& E, negedge D, `FD7HS_D_CP_SETUP_negedge_posedge, `FD7HS_D_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP, posedge E, `FD7HS_E_CP_SETUP_posedge_posedge, `FD7HS_E_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP, negedge E, `FD7HS_E_CP_SETUP_negedge_posedge, `FD7HS_E_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD7HS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7HS_CP_PWH, 0, Notifier);
 
   endspecify
`endif
 
endmodule // FD7HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:57 and Version :1.1 //
 
//  START 
// CELL FD7HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD7HSP_CP_R_QN_F 0.1
`define FD7HSP_CP_R_QN_R 0.1
`define FD7HSP_CP_R_Q_R 0.1
`define FD7HSP_CP_R_Q_F 0.1
`define FD7HSP_CP_PWH 0.1
`define FD7HSP_CP_PWL 0.1
`define FD7HSP_E_CP_SETUP_posedge_posedge 0.1
`define FD7HSP_E_CP_SETUP_negedge_posedge 0.1
`define FD7HSP_E_CP_HOLD_posedge_posedge 0.1
`define FD7HSP_E_CP_HOLD_negedge_posedge 0.1
`define FD7HSP_D_CP_SETUP_posedge_posedge 0.1
`define FD7HSP_D_CP_SETUP_negedge_posedge 0.1
`define FD7HSP_D_CP_HOLD_posedge_posedge 0.1
`define FD7HSP_D_CP_HOLD_negedge_posedge 0.1
 
module FD7HSP (Q, QN, D, E, CP);
 
   output Q;
   output QN;
   input D;
   input E;
   input CP;
 
 
   reg Notifier;
 
   U_MUX2  u0 (Mux21IQDE_, IQ, D, E);
 
   U_FD_P_NOTI u2 (   // Verilog Seq UDP
     IQ, Mux21IQDE_, CP, Notifier);
 
   buf  u3 (Q, IQ);
   not  u4 (QN, IQ);
 
 
 
`ifdef functional
`else
   specify
 
      (posedge CP => (Q +: D)) = (`FD7HSP_CP_R_Q_R, `FD7HSP_CP_R_Q_F);
      (posedge CP => (QN -: D)) = (`FD7HSP_CP_R_QN_R, `FD7HSP_CP_R_QN_F);
 
	$setuphold(posedge CP &&& E, posedge D, `FD7HSP_D_CP_SETUP_posedge_posedge, `FD7HSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& E, negedge D, `FD7HSP_D_CP_SETUP_negedge_posedge, `FD7HSP_D_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP, posedge E, `FD7HSP_E_CP_SETUP_posedge_posedge, `FD7HSP_E_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP, negedge E, `FD7HSP_E_CP_SETUP_negedge_posedge, `FD7HSP_E_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD7HSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7HSP_CP_PWH, 0, Notifier);
 
   endspecify
`endif
 
endmodule // FD7HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:57 and Version :1.1 //
 
//  START 
// CELL FD7SHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD7SHS_CP_R_QN_F 0.1
`define FD7SHS_CP_R_QN_R 0.1
`define FD7SHS_CP_R_Q_R 0.1
`define FD7SHS_CP_R_Q_F 0.1
`define FD7SHS_CP_PWH 0.1
`define FD7SHS_CP_PWL 0.1
`define FD7SHS_TE_CP_SETUP_posedge_posedge 0.1
`define FD7SHS_TE_CP_SETUP_negedge_posedge 0.1
`define FD7SHS_TE_CP_HOLD_posedge_posedge 0.1
`define FD7SHS_TE_CP_HOLD_negedge_posedge 0.1
`define FD7SHS_TI_CP_SETUP_posedge_posedge 0.1
`define FD7SHS_TI_CP_SETUP_negedge_posedge 0.1
`define FD7SHS_TI_CP_HOLD_posedge_posedge 0.1
`define FD7SHS_TI_CP_HOLD_negedge_posedge 0.1
`define FD7SHS_E_CP_SETUP_posedge_posedge 0.1
`define FD7SHS_E_CP_SETUP_negedge_posedge 0.1
`define FD7SHS_E_CP_HOLD_posedge_posedge 0.1
`define FD7SHS_E_CP_HOLD_negedge_posedge 0.1
`define FD7SHS_D_CP_SETUP_posedge_posedge 0.1
`define FD7SHS_D_CP_SETUP_negedge_posedge 0.1
`define FD7SHS_D_CP_HOLD_posedge_posedge 0.1
`define FD7SHS_D_CP_HOLD_negedge_posedge 0.1
 
module FD7SHS (Q, QN, D, E, CP, TI, TE);
 
   output Q;
   output QN;
   input CP;
   input TE;
   input TI;
   input E;
   input D;
 
 
   reg Notifier;
 
   U_MUX2  u0 (Mux21IQDE_, IQ, D, E);
   U_MUX2  u1 (Mux21Mux21IQDE_TITE_, Mux21IQDE_, TI, TE);
 
   U_FD_P_NOTI u2 (   // Verilog Seq UDP
     IQ, Mux21Mux21IQDE_TITE_, CP, Notifier);
 
   buf  u3 (Q, IQ);
   not  u4 (QN, IQ);
 
 
 
`ifdef functional
`else
   and  (DE_, D, E);
   and  (QE_, Q, E_);
    or  (DEor_, DE_, QE_);
   not  (E_, E);

   xor  (D_orTI, DEor_, TI);
   not  (TEX, TE);
   and  (AndTEXE_, TEX, E);
   specify
`ifdef verifault
 
      if(!IQ && !E && TI) (posedge CP => (Q +: TE)) = (`FD7SHS_CP_R_Q_R, `FD7SHS_CP_R_Q_F);
      if(!D && E && TI) (posedge CP => (Q +: TE)) = (`FD7SHS_CP_R_Q_R, `FD7SHS_CP_R_Q_F);
      if(!TI && E && D) (posedge CP => (Q -: TE)) = (`FD7SHS_CP_R_Q_R, `FD7SHS_CP_R_Q_F);
      if(!TI && !E && IQ) (posedge CP => (Q -: TE)) = (`FD7SHS_CP_R_Q_R, `FD7SHS_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD7SHS_CP_R_Q_R, `FD7SHS_CP_R_Q_F);
      if(!IQ && !TE && D) (posedge CP => (Q +: E)) = (`FD7SHS_CP_R_Q_R, `FD7SHS_CP_R_Q_F);
      if(!D && !TE && IQ) (posedge CP => (Q -: E)) = (`FD7SHS_CP_R_Q_R, `FD7SHS_CP_R_Q_F);
      if(!TE && E) (posedge CP => (Q +: D)) = (`FD7SHS_CP_R_Q_R, `FD7SHS_CP_R_Q_F);
      if(!IQ && !E && TI) (posedge CP => (QN -: TE)) = (`FD7SHS_CP_R_QN_R, `FD7SHS_CP_R_QN_F);
      if(!D && E && TI) (posedge CP => (QN -: TE)) = (`FD7SHS_CP_R_QN_R, `FD7SHS_CP_R_QN_F);
      if(!TI && E && D) (posedge CP => (QN +: TE)) = (`FD7SHS_CP_R_QN_R, `FD7SHS_CP_R_QN_F);
      if(!TI && !E && IQ) (posedge CP => (QN +: TE)) = (`FD7SHS_CP_R_QN_R, `FD7SHS_CP_R_QN_F);
      if(TE) (posedge CP => (QN -: TI)) = (`FD7SHS_CP_R_QN_R, `FD7SHS_CP_R_QN_F);
      if(!IQ && !TE && D) (posedge CP => (QN -: E)) = (`FD7SHS_CP_R_QN_R, `FD7SHS_CP_R_QN_F);
      if(!D && !TE && IQ) (posedge CP => (QN +: E)) = (`FD7SHS_CP_R_QN_R, `FD7SHS_CP_R_QN_F);
      if(!TE && E) (posedge CP => (QN -: D)) = (`FD7SHS_CP_R_QN_R, `FD7SHS_CP_R_QN_F);
 
	$setuphold(posedge CP &&& AndTEXE_, posedge D, `FD7SHS_D_CP_SETUP_posedge_posedge, `FD7SHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndTEXE_, negedge D, `FD7SHS_D_CP_SETUP_negedge_posedge, `FD7SHS_D_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TEX, posedge E, `FD7SHS_E_CP_SETUP_posedge_posedge, `FD7SHS_E_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TEX, negedge E, `FD7SHS_E_CP_SETUP_negedge_posedge, `FD7SHS_E_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FD7SHS_TI_CP_SETUP_posedge_posedge, `FD7SHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FD7SHS_TI_CP_SETUP_negedge_posedge, `FD7SHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& D_orTI, posedge TE, `FD7SHS_TE_CP_SETUP_posedge_posedge, `FD7SHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& D_orTI, negedge TE, `FD7SHS_TE_CP_SETUP_negedge_posedge, `FD7SHS_TE_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD7SHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7SHS_CP_PWH, 0, Notifier);
`else
 
      (posedge CP => (Q +: Mux21Mux21IQDE_TITE_)) = (`FD7SHS_CP_R_Q_R, `FD7SHS_CP_R_Q_F);
      (posedge CP => (QN -: Mux21Mux21IQDE_TITE_)) = (`FD7SHS_CP_R_QN_R, `FD7SHS_CP_R_QN_F);
 
        $setuphold(posedge CP &&& AndTEXE_, posedge D, `FD7SHS_D_CP_SETUP_posedge_posedge, `FD7SHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndTEXE_, negedge D, `FD7SHS_D_CP_SETUP_negedge_posedge, `FD7SHS_D_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge E, `FD7SHS_E_CP_SETUP_posedge_posedge, `FD7SHS_E_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge E, `FD7SHS_E_CP_SETUP_negedge_posedge, `FD7SHS_E_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD7SHS_TI_CP_SETUP_posedge_posedge, `FD7SHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD7SHS_TI_CP_SETUP_negedge_posedge, `FD7SHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& D_orTI, posedge TE, `FD7SHS_TE_CP_SETUP_posedge_posedge, `FD7SHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& D_orTI, negedge TE, `FD7SHS_TE_CP_SETUP_negedge_posedge, `FD7SHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD7SHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7SHS_CP_PWH, 0, Notifier);
`endif 
   endspecify
`endif
 
endmodule // FD7SHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:57 and Version :1.1 //
 
//  START 
// CELL FD7SHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD7SHSP_CP_R_QN_F 0.1
`define FD7SHSP_CP_R_QN_R 0.1
`define FD7SHSP_CP_R_Q_R 0.1
`define FD7SHSP_CP_R_Q_F 0.1
`define FD7SHSP_CP_PWH 0.1
`define FD7SHSP_CP_PWL 0.1
`define FD7SHSP_TE_CP_SETUP_posedge_posedge 0.1
`define FD7SHSP_TE_CP_SETUP_negedge_posedge 0.1
`define FD7SHSP_TE_CP_HOLD_posedge_posedge 0.1
`define FD7SHSP_TE_CP_HOLD_negedge_posedge 0.1
`define FD7SHSP_TI_CP_SETUP_posedge_posedge 0.1
`define FD7SHSP_TI_CP_SETUP_negedge_posedge 0.1
`define FD7SHSP_TI_CP_HOLD_posedge_posedge 0.1
`define FD7SHSP_TI_CP_HOLD_negedge_posedge 0.1
`define FD7SHSP_E_CP_SETUP_posedge_posedge 0.1
`define FD7SHSP_E_CP_SETUP_negedge_posedge 0.1
`define FD7SHSP_E_CP_HOLD_posedge_posedge 0.1
`define FD7SHSP_E_CP_HOLD_negedge_posedge 0.1
`define FD7SHSP_D_CP_SETUP_posedge_posedge 0.1
`define FD7SHSP_D_CP_SETUP_negedge_posedge 0.1
`define FD7SHSP_D_CP_HOLD_posedge_posedge 0.1
`define FD7SHSP_D_CP_HOLD_negedge_posedge 0.1
 
module FD7SHSP (Q, QN, D, E, CP, TI, TE);
 
   output Q;
   output QN;
   input CP;
   input TE;
   input TI;
   input E;
   input D;
 
 
   reg Notifier;
 
   U_MUX2  u0 (Mux21IQDE_, IQ, D, E);
   U_MUX2  u1 (Mux21Mux21IQDE_TITE_, Mux21IQDE_, TI, TE);
 
   U_FD_P_NOTI u2 (   // Verilog Seq UDP
     IQ, Mux21Mux21IQDE_TITE_, CP, Notifier);
 
   buf  u3 (Q, IQ);
   not  u4 (QN, IQ);
 
 
 
`ifdef functional
`else
   and  (DE_, D, E);
   and  (QE_, Q, E_);
    or  (DEor_, DE_, QE_);
   not  (E_, E);

   xor  (D_orTI, DEor_, TI);
   not  (TEX, TE);
   and  (AndTEXE_, TEX, E);
   specify
`ifdef verifault
 
      if(!IQ && !E && TI) (posedge CP => (Q +: TE)) = (`FD7SHSP_CP_R_Q_R, `FD7SHSP_CP_R_Q_F);
      if(!D && E && TI) (posedge CP => (Q +: TE)) = (`FD7SHSP_CP_R_Q_R, `FD7SHSP_CP_R_Q_F);
      if(!TI && E && D) (posedge CP => (Q -: TE)) = (`FD7SHSP_CP_R_Q_R, `FD7SHSP_CP_R_Q_F);
      if(!TI && !E && IQ) (posedge CP => (Q -: TE)) = (`FD7SHSP_CP_R_Q_R, `FD7SHSP_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD7SHSP_CP_R_Q_R, `FD7SHSP_CP_R_Q_F);
      if(!IQ && !TE && D) (posedge CP => (Q +: E)) = (`FD7SHSP_CP_R_Q_R, `FD7SHSP_CP_R_Q_F);
      if(!D && !TE && IQ) (posedge CP => (Q -: E)) = (`FD7SHSP_CP_R_Q_R, `FD7SHSP_CP_R_Q_F);
      if(!TE && E) (posedge CP => (Q +: D)) = (`FD7SHSP_CP_R_Q_R, `FD7SHSP_CP_R_Q_F);
      if(!IQ && !E && TI) (posedge CP => (QN -: TE)) = (`FD7SHSP_CP_R_QN_R, `FD7SHSP_CP_R_QN_F);
      if(!D && E && TI) (posedge CP => (QN -: TE)) = (`FD7SHSP_CP_R_QN_R, `FD7SHSP_CP_R_QN_F);
      if(!TI && E && D) (posedge CP => (QN +: TE)) = (`FD7SHSP_CP_R_QN_R, `FD7SHSP_CP_R_QN_F);
      if(!TI && !E && IQ) (posedge CP => (QN +: TE)) = (`FD7SHSP_CP_R_QN_R, `FD7SHSP_CP_R_QN_F);
      if(TE) (posedge CP => (QN -: TI)) = (`FD7SHSP_CP_R_QN_R, `FD7SHSP_CP_R_QN_F);
      if(!IQ && !TE && D) (posedge CP => (QN -: E)) = (`FD7SHSP_CP_R_QN_R, `FD7SHSP_CP_R_QN_F);
      if(!D && !TE && IQ) (posedge CP => (QN +: E)) = (`FD7SHSP_CP_R_QN_R, `FD7SHSP_CP_R_QN_F);
      if(!TE && E) (posedge CP => (QN -: D)) = (`FD7SHSP_CP_R_QN_R, `FD7SHSP_CP_R_QN_F);
 
	$setuphold(posedge CP &&& AndTEXE_, posedge D, `FD7SHSP_D_CP_SETUP_posedge_posedge, `FD7SHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndTEXE_, negedge D, `FD7SHSP_D_CP_SETUP_negedge_posedge, `FD7SHSP_D_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TEX, posedge E, `FD7SHSP_E_CP_SETUP_posedge_posedge, `FD7SHSP_E_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TEX, negedge E, `FD7SHSP_E_CP_SETUP_negedge_posedge, `FD7SHSP_E_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FD7SHSP_TI_CP_SETUP_posedge_posedge, `FD7SHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FD7SHSP_TI_CP_SETUP_negedge_posedge, `FD7SHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& D_orTI, posedge TE, `FD7SHSP_TE_CP_SETUP_posedge_posedge, `FD7SHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& D_orTI, negedge TE, `FD7SHSP_TE_CP_SETUP_negedge_posedge, `FD7SHSP_TE_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD7SHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7SHSP_CP_PWH, 0, Notifier);
`else
 
      (posedge CP => (Q +: Mux21Mux21IQDE_TITE_)) = (`FD7SHSP_CP_R_Q_R, `FD7SHSP_CP_R_Q_F);
      (posedge CP => (QN -: Mux21Mux21IQDE_TITE_)) = (`FD7SHSP_CP_R_QN_R, `FD7SHSP_CP_R_QN_F);
 
        $setuphold(posedge CP &&& AndTEXE_, posedge D, `FD7SHSP_D_CP_SETUP_posedge_posedge, `FD7SHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndTEXE_, negedge D, `FD7SHSP_D_CP_SETUP_negedge_posedge, `FD7SHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge E, `FD7SHSP_E_CP_SETUP_posedge_posedge, `FD7SHSP_E_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge E, `FD7SHSP_E_CP_SETUP_negedge_posedge, `FD7SHSP_E_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD7SHSP_TI_CP_SETUP_posedge_posedge, `FD7SHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD7SHSP_TI_CP_SETUP_negedge_posedge, `FD7SHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& D_orTI, posedge TE, `FD7SHSP_TE_CP_SETUP_posedge_posedge, `FD7SHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& D_orTI, negedge TE, `FD7SHSP_TE_CP_SETUP_negedge_posedge, `FD7SHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD7SHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7SHSP_CP_PWH, 0, Notifier);
`endif 
   endspecify
`endif
 
endmodule // FD7SHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:57 and Version :1.1 //
 
//  START 
// CELL FD7SQHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD7SQHS_CP_R_Q_R 0.1
`define FD7SQHS_CP_R_Q_F 0.1
`define FD7SQHS_CP_PWH 0.1
`define FD7SQHS_CP_PWL 0.1
`define FD7SQHS_TE_CP_SETUP_posedge_posedge 0.1
`define FD7SQHS_TE_CP_SETUP_negedge_posedge 0.1
`define FD7SQHS_TE_CP_HOLD_posedge_posedge 0.1
`define FD7SQHS_TE_CP_HOLD_negedge_posedge 0.1
`define FD7SQHS_TI_CP_SETUP_posedge_posedge 0.1
`define FD7SQHS_TI_CP_SETUP_negedge_posedge 0.1
`define FD7SQHS_TI_CP_HOLD_posedge_posedge 0.1
`define FD7SQHS_TI_CP_HOLD_negedge_posedge 0.1
`define FD7SQHS_E_CP_SETUP_posedge_posedge 0.1
`define FD7SQHS_E_CP_SETUP_negedge_posedge 0.1
`define FD7SQHS_E_CP_HOLD_posedge_posedge 0.1
`define FD7SQHS_E_CP_HOLD_negedge_posedge 0.1
`define FD7SQHS_D_CP_SETUP_posedge_posedge 0.1
`define FD7SQHS_D_CP_SETUP_negedge_posedge 0.1
`define FD7SQHS_D_CP_HOLD_posedge_posedge 0.1
`define FD7SQHS_D_CP_HOLD_negedge_posedge 0.1
 
module FD7SQHS (Q, D, E, CP, TI, TE);
 
   output Q;
   input CP;
   input TE;
   input TI;
   input E;
   input D;
 
 
   reg Notifier;
 
   U_MUX2  u0 (Mux21IQDE_, IQ, D, E);
   U_MUX2  u1 (Mux21Mux21IQDE_TITE_, Mux21IQDE_, TI, TE);
 
   U_FD_P_NOTI u2 (   // Verilog Seq UDP
      IQ, Mux21Mux21IQDE_TITE_, CP, Notifier);
 
   buf  u3 (Q, IQ);
 
 
 
`ifdef functional
`else
   and  (DE_, D, E);
   and  (QE_, Q, E_);
    or  (DEor_, DE_, QE_);
   not  (E_, E);

   xor  (D_orTI, DEor_, TI);
   not  (TEX, TE);
   and  (AndTEXE_, TEX, E);
   specify
`ifdef verifault 
      if(!IQ && !E && TI) (posedge CP => (Q +: TE)) = (`FD7SQHS_CP_R_Q_R, `FD7SQHS_CP_R_Q_F);
      if(!D && E && TI) (posedge CP => (Q +: TE)) = (`FD7SQHS_CP_R_Q_R, `FD7SQHS_CP_R_Q_F);
      if(!TI && E && D) (posedge CP => (Q -: TE)) = (`FD7SQHS_CP_R_Q_R, `FD7SQHS_CP_R_Q_F);
      if(!TI && !E && IQ) (posedge CP => (Q -: TE)) = (`FD7SQHS_CP_R_Q_R, `FD7SQHS_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD7SQHS_CP_R_Q_R, `FD7SQHS_CP_R_Q_F);
      if(!IQ && !TE && D) (posedge CP => (Q +: E)) = (`FD7SQHS_CP_R_Q_R, `FD7SQHS_CP_R_Q_F);
      if(!D && !TE && IQ) (posedge CP => (Q -: E)) = (`FD7SQHS_CP_R_Q_R, `FD7SQHS_CP_R_Q_F);
      if(!TE && E) (posedge CP => (Q +: D)) = (`FD7SQHS_CP_R_Q_R, `FD7SQHS_CP_R_Q_F);
 
	$setuphold(posedge CP &&& AndTEXE_, posedge D, `FD7SQHS_D_CP_SETUP_posedge_posedge, `FD7SQHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndTEXE_, negedge D, `FD7SQHS_D_CP_SETUP_negedge_posedge, `FD7SQHS_D_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TEX, posedge E, `FD7SQHS_E_CP_SETUP_posedge_posedge, `FD7SQHS_E_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TEX, negedge E, `FD7SQHS_E_CP_SETUP_negedge_posedge, `FD7SQHS_E_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FD7SQHS_TI_CP_SETUP_posedge_posedge, `FD7SQHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FD7SQHS_TI_CP_SETUP_negedge_posedge, `FD7SQHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& D_orTI, posedge TE, `FD7SQHS_TE_CP_SETUP_posedge_posedge, `FD7SQHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& D_orTI, negedge TE, `FD7SQHS_TE_CP_SETUP_negedge_posedge, `FD7SQHS_TE_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD7SQHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7SQHS_CP_PWH, 0, Notifier);
`else
      (posedge CP => (Q +: Mux21Mux21IQDE_TITE_)) = (`FD7SQHS_CP_R_Q_R, `FD7SQHS_CP_R_Q_F);
 
        $setuphold(posedge CP &&& AndTEXE_, posedge D, `FD7SQHS_D_CP_SETUP_posedge_posedge, `FD7SQHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndTEXE_, negedge D, `FD7SQHS_D_CP_SETUP_negedge_posedge, `FD7SQHS_D_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge E, `FD7SQHS_E_CP_SETUP_posedge_posedge, `FD7SQHS_E_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge E, `FD7SQHS_E_CP_SETUP_negedge_posedge, `FD7SQHS_E_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD7SQHS_TI_CP_SETUP_posedge_posedge, `FD7SQHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD7SQHS_TI_CP_SETUP_negedge_posedge, `FD7SQHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& D_orTI, posedge TE, `FD7SQHS_TE_CP_SETUP_posedge_posedge, `FD7SQHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& D_orTI, negedge TE, `FD7SQHS_TE_CP_SETUP_negedge_posedge, `FD7SQHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD7SQHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7SQHS_CP_PWH, 0, Notifier);
 `endif 
   endspecify
`endif
 
 
endmodule // FD7SQHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:01 and Version :1.1 //
 
//  START 
// CELL FD7SQHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD7SQHSP_CP_R_Q_R 0.1
`define FD7SQHSP_CP_R_Q_F 0.1
`define FD7SQHSP_CP_PWH 0.1
`define FD7SQHSP_CP_PWL 0.1
`define FD7SQHSP_TE_CP_SETUP_posedge_posedge 0.1
`define FD7SQHSP_TE_CP_SETUP_negedge_posedge 0.1
`define FD7SQHSP_TE_CP_HOLD_posedge_posedge 0.1
`define FD7SQHSP_TE_CP_HOLD_negedge_posedge 0.1
`define FD7SQHSP_TI_CP_SETUP_posedge_posedge 0.1
`define FD7SQHSP_TI_CP_SETUP_negedge_posedge 0.1
`define FD7SQHSP_TI_CP_HOLD_posedge_posedge 0.1
`define FD7SQHSP_TI_CP_HOLD_negedge_posedge 0.1
`define FD7SQHSP_E_CP_SETUP_posedge_posedge 0.1
`define FD7SQHSP_E_CP_SETUP_negedge_posedge 0.1
`define FD7SQHSP_E_CP_HOLD_posedge_posedge 0.1
`define FD7SQHSP_E_CP_HOLD_negedge_posedge 0.1
`define FD7SQHSP_D_CP_SETUP_posedge_posedge 0.1
`define FD7SQHSP_D_CP_SETUP_negedge_posedge 0.1
`define FD7SQHSP_D_CP_HOLD_posedge_posedge 0.1
`define FD7SQHSP_D_CP_HOLD_negedge_posedge 0.1
 
module FD7SQHSP (Q, D, E, CP, TI, TE);
 
   output Q;
   input CP;
   input TE;
   input TI;
   input E;
   input D;
 
 
   reg Notifier;
 
   U_MUX2  u0 (Mux21IQDE_, IQ, D, E);
   U_MUX2  u1 (Mux21Mux21IQDE_TITE_, Mux21IQDE_, TI, TE);
 
   U_FD_P_NOTI u2 (   // Verilog Seq UDP
      IQ, Mux21Mux21IQDE_TITE_, CP, Notifier);
 
   buf  u3 (Q, IQ);
 
 
 
`ifdef functional
`else
   and  (DE_, D, E);
   and  (QE_, Q, E_);
    or  (DEor_, DE_, QE_);
   not  (E_, E);

   xor  (D_orTI, DEor_, TI);
   not  (TEX, TE);
   and  (AndTEXE_, TEX, E);
   specify
`ifdef verifault 
      if(!IQ && !E && TI) (posedge CP => (Q +: TE)) = (`FD7SQHSP_CP_R_Q_R, `FD7SQHSP_CP_R_Q_F);
      if(!D && E && TI) (posedge CP => (Q +: TE)) = (`FD7SQHSP_CP_R_Q_R, `FD7SQHSP_CP_R_Q_F);
      if(!TI && E && D) (posedge CP => (Q -: TE)) = (`FD7SQHSP_CP_R_Q_R, `FD7SQHSP_CP_R_Q_F);
      if(!TI && !E && IQ) (posedge CP => (Q -: TE)) = (`FD7SQHSP_CP_R_Q_R, `FD7SQHSP_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD7SQHSP_CP_R_Q_R, `FD7SQHSP_CP_R_Q_F);
      if(!IQ && !TE && D) (posedge CP => (Q +: E)) = (`FD7SQHSP_CP_R_Q_R, `FD7SQHSP_CP_R_Q_F);
      if(!D && !TE && IQ) (posedge CP => (Q -: E)) = (`FD7SQHSP_CP_R_Q_R, `FD7SQHSP_CP_R_Q_F);
      if(!TE && E) (posedge CP => (Q +: D)) = (`FD7SQHSP_CP_R_Q_R, `FD7SQHSP_CP_R_Q_F);
 
	$setuphold(posedge CP &&& AndTEXE_, posedge D, `FD7SQHSP_D_CP_SETUP_posedge_posedge, `FD7SQHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndTEXE_, negedge D, `FD7SQHSP_D_CP_SETUP_negedge_posedge, `FD7SQHSP_D_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TEX, posedge E, `FD7SQHSP_E_CP_SETUP_posedge_posedge, `FD7SQHSP_E_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TEX, negedge E, `FD7SQHSP_E_CP_SETUP_negedge_posedge, `FD7SQHSP_E_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FD7SQHSP_TI_CP_SETUP_posedge_posedge, `FD7SQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FD7SQHSP_TI_CP_SETUP_negedge_posedge, `FD7SQHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& D_orTI, posedge TE, `FD7SQHSP_TE_CP_SETUP_posedge_posedge, `FD7SQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& D_orTI, negedge TE, `FD7SQHSP_TE_CP_SETUP_negedge_posedge, `FD7SQHSP_TE_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD7SQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7SQHSP_CP_PWH, 0, Notifier);
`else
      (posedge CP => (Q +: Mux21Mux21IQDE_TITE_)) = (`FD7SQHSP_CP_R_Q_R, `FD7SQHSP_CP_R_Q_F);
 
        $setuphold(posedge CP &&& AndTEXE_, posedge D, `FD7SQHSP_D_CP_SETUP_posedge_posedge, `FD7SQHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndTEXE_, negedge D, `FD7SQHSP_D_CP_SETUP_negedge_posedge, `FD7SQHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge E, `FD7SQHSP_E_CP_SETUP_posedge_posedge, `FD7SQHSP_E_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge E, `FD7SQHSP_E_CP_SETUP_negedge_posedge, `FD7SQHSP_E_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD7SQHSP_TI_CP_SETUP_posedge_posedge, `FD7SQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD7SQHSP_TI_CP_SETUP_negedge_posedge, `FD7SQHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& D_orTI, posedge TE, `FD7SQHSP_TE_CP_SETUP_posedge_posedge, `FD7SQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& D_orTI, negedge TE, `FD7SQHSP_TE_CP_SETUP_negedge_posedge, `FD7SQHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD7SQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7SQHSP_CP_PWH, 0, Notifier);
 `endif 
   endspecify
`endif
 
 
endmodule // FD7SQHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:01 and Version :1.1 //
 
//  START 
// CELL FD7SQHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD7SQHSX4_CP_R_Q_R 0.1
`define FD7SQHSX4_CP_R_Q_F 0.1
`define FD7SQHSX4_CP_PWH 0.1
`define FD7SQHSX4_CP_PWL 0.1
`define FD7SQHSX4_TE_CP_SETUP_posedge_posedge 0.1
`define FD7SQHSX4_TE_CP_SETUP_negedge_posedge 0.1
`define FD7SQHSX4_TE_CP_HOLD_posedge_posedge 0.1
`define FD7SQHSX4_TE_CP_HOLD_negedge_posedge 0.1
`define FD7SQHSX4_TI_CP_SETUP_posedge_posedge 0.1
`define FD7SQHSX4_TI_CP_SETUP_negedge_posedge 0.1
`define FD7SQHSX4_TI_CP_HOLD_posedge_posedge 0.1
`define FD7SQHSX4_TI_CP_HOLD_negedge_posedge 0.1
`define FD7SQHSX4_E_CP_SETUP_posedge_posedge 0.1
`define FD7SQHSX4_E_CP_SETUP_negedge_posedge 0.1
`define FD7SQHSX4_E_CP_HOLD_posedge_posedge 0.1
`define FD7SQHSX4_E_CP_HOLD_negedge_posedge 0.1
`define FD7SQHSX4_D_CP_SETUP_posedge_posedge 0.1
`define FD7SQHSX4_D_CP_SETUP_negedge_posedge 0.1
`define FD7SQHSX4_D_CP_HOLD_posedge_posedge 0.1
`define FD7SQHSX4_D_CP_HOLD_negedge_posedge 0.1
 
module FD7SQHSX4 (Q, D, E, CP, TI, TE);
 
   output Q;
   input CP;
   input TE;
   input TI;
   input E;
   input D;
 
 
   reg Notifier;
 
   U_MUX2  u0 (Mux21IQDE_, IQ, D, E);
   U_MUX2  u1 (Mux21Mux21IQDE_TITE_, Mux21IQDE_, TI, TE);
 
   U_FD_P_NOTI u2 (   // Verilog Seq UDP
      IQ, Mux21Mux21IQDE_TITE_, CP, Notifier);
 
   buf  u3 (Q, IQ);
 
 
 
`ifdef functional
`else
   and  (DE_, D, E);
   and  (QE_, Q, E_);
    or  (DEor_, DE_, QE_);
   not  (E_, E);

   xor  (D_orTI, DEor_, TI);
   not  (TEX, TE);
   and  (AndTEXE_, TEX, E);
   specify
`ifdef verifault 
      if(!IQ && !E && TI) (posedge CP => (Q +: TE)) = (`FD7SQHSX4_CP_R_Q_R, `FD7SQHSX4_CP_R_Q_F);
      if(!D && E && TI) (posedge CP => (Q +: TE)) = (`FD7SQHSX4_CP_R_Q_R, `FD7SQHSX4_CP_R_Q_F);
      if(!TI && E && D) (posedge CP => (Q -: TE)) = (`FD7SQHSX4_CP_R_Q_R, `FD7SQHSX4_CP_R_Q_F);
      if(!TI && !E && IQ) (posedge CP => (Q -: TE)) = (`FD7SQHSX4_CP_R_Q_R, `FD7SQHSX4_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD7SQHSX4_CP_R_Q_R, `FD7SQHSX4_CP_R_Q_F);
      if(!IQ && !TE && D) (posedge CP => (Q +: E)) = (`FD7SQHSX4_CP_R_Q_R, `FD7SQHSX4_CP_R_Q_F);
      if(!D && !TE && IQ) (posedge CP => (Q -: E)) = (`FD7SQHSX4_CP_R_Q_R, `FD7SQHSX4_CP_R_Q_F);
      if(!TE && E) (posedge CP => (Q +: D)) = (`FD7SQHSX4_CP_R_Q_R, `FD7SQHSX4_CP_R_Q_F);
 
	$setuphold(posedge CP &&& AndTEXE_, posedge D, `FD7SQHSX4_D_CP_SETUP_posedge_posedge, `FD7SQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndTEXE_, negedge D, `FD7SQHSX4_D_CP_SETUP_negedge_posedge, `FD7SQHSX4_D_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TEX, posedge E, `FD7SQHSX4_E_CP_SETUP_posedge_posedge, `FD7SQHSX4_E_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TEX, negedge E, `FD7SQHSX4_E_CP_SETUP_negedge_posedge, `FD7SQHSX4_E_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FD7SQHSX4_TI_CP_SETUP_posedge_posedge, `FD7SQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FD7SQHSX4_TI_CP_SETUP_negedge_posedge, `FD7SQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& D_orTI, posedge TE, `FD7SQHSX4_TE_CP_SETUP_posedge_posedge, `FD7SQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& D_orTI, negedge TE, `FD7SQHSX4_TE_CP_SETUP_negedge_posedge, `FD7SQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD7SQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7SQHSX4_CP_PWH, 0, Notifier);
`else
      (posedge CP => (Q +: Mux21Mux21IQDE_TITE_)) = (`FD7SQHSX4_CP_R_Q_R, `FD7SQHSX4_CP_R_Q_F);
 
        $setuphold(posedge CP &&& AndTEXE_, posedge D, `FD7SQHSX4_D_CP_SETUP_posedge_posedge, `FD7SQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndTEXE_, negedge D, `FD7SQHSX4_D_CP_SETUP_negedge_posedge, `FD7SQHSX4_D_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge E, `FD7SQHSX4_E_CP_SETUP_posedge_posedge, `FD7SQHSX4_E_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge E, `FD7SQHSX4_E_CP_SETUP_negedge_posedge, `FD7SQHSX4_E_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD7SQHSX4_TI_CP_SETUP_posedge_posedge, `FD7SQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD7SQHSX4_TI_CP_SETUP_negedge_posedge, `FD7SQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& D_orTI, posedge TE, `FD7SQHSX4_TE_CP_SETUP_posedge_posedge, `FD7SQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& D_orTI, negedge TE, `FD7SQHSX4_TE_CP_SETUP_negedge_posedge, `FD7SQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD7SQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7SQHSX4_CP_PWH, 0, Notifier);
 `endif 
   endspecify
`endif
 
 
endmodule // FD7SQHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:01 and Version :1.1 //
 
//  START 
// CELL FD7THS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD7THS_CP_R_QN_F 0.1
`define FD7THS_CP_R_QN_R 0.1
`define FD7THS_CP_R_Q_R 0.1
`define FD7THS_CP_R_Q_F 0.1
`define FD7THS_CP_R_SO_R 0.1
`define FD7THS_CP_R_SO_F 0.1
`define FD7THS_CP_PWH 0.1
`define FD7THS_CP_PWL 0.1
`define FD7THS_TE_CP_SETUP_posedge_posedge 0.1
`define FD7THS_TE_CP_SETUP_negedge_posedge 0.1
`define FD7THS_TE_CP_HOLD_posedge_posedge 0.1
`define FD7THS_TE_CP_HOLD_negedge_posedge 0.1
`define FD7THS_TI_CP_SETUP_posedge_posedge 0.1
`define FD7THS_TI_CP_SETUP_negedge_posedge 0.1
`define FD7THS_TI_CP_HOLD_posedge_posedge 0.1
`define FD7THS_TI_CP_HOLD_negedge_posedge 0.1
`define FD7THS_E_CP_SETUP_posedge_posedge 0.1
`define FD7THS_E_CP_SETUP_negedge_posedge 0.1
`define FD7THS_E_CP_HOLD_posedge_posedge 0.1
`define FD7THS_E_CP_HOLD_negedge_posedge 0.1
`define FD7THS_D_CP_SETUP_posedge_posedge 0.1
`define FD7THS_D_CP_SETUP_negedge_posedge 0.1
`define FD7THS_D_CP_HOLD_posedge_posedge 0.1
`define FD7THS_D_CP_HOLD_negedge_posedge 0.1
 
module FD7THS (Q, QN, SO, D, E, CP, TI, TE);
 
   output Q;
   output QN;
   output SO;
   input CP;
   input TE;
   input TI;
   input E;
   input D;
 
 
   reg Notifier;
 
   U_MUX2  u0 (Mux21IQDE_, IQ, D, E);
   U_MUX2  u1 (Mux21Mux21IQDE_TITE_, Mux21IQDE_, TI, TE);
 
   U_FD_P_NOTI u2 (   // Verilog Seq UDP
     IQ, Mux21Mux21IQDE_TITE_, CP, Notifier);
 
   buf  u3 (Q, IQ);
   not  u4 (QN, IQ);
   buf  u5 (SO, IQ);
 
 
 
`ifdef functional
`else
   and  (DE_, D, E);
   and  (QE_, Q, E_);
    or  (DEor_, DE_, QE_);
   not  (E_, E);

   xor  (D_orTI, DEor_, TI);
   not  (TEX, TE);
   and  (AndTEXE_, TEX, E);
   specify
`ifdef verifault
 
      if(!IQ && !E && TI) (posedge CP => (Q +: TE)) = (`FD7THS_CP_R_Q_R, `FD7THS_CP_R_Q_F);
      if(!D && E && TI) (posedge CP => (Q +: TE)) = (`FD7THS_CP_R_Q_R, `FD7THS_CP_R_Q_F);
      if(!TI && E && D) (posedge CP => (Q -: TE)) = (`FD7THS_CP_R_Q_R, `FD7THS_CP_R_Q_F);
      if(!TI && !E && IQ) (posedge CP => (Q -: TE)) = (`FD7THS_CP_R_Q_R, `FD7THS_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD7THS_CP_R_Q_R, `FD7THS_CP_R_Q_F);
      if(!IQ && !TE && D) (posedge CP => (Q +: E)) = (`FD7THS_CP_R_Q_R, `FD7THS_CP_R_Q_F);
      if(!D && !TE && IQ) (posedge CP => (Q -: E)) = (`FD7THS_CP_R_Q_R, `FD7THS_CP_R_Q_F);
      if(!TE && E) (posedge CP => (Q +: D)) = (`FD7THS_CP_R_Q_R, `FD7THS_CP_R_Q_F);
      if(!IQ && !E && TI) (posedge CP => (QN -: TE)) = (`FD7THS_CP_R_QN_R, `FD7THS_CP_R_QN_F);
      if(!D && E && TI) (posedge CP => (QN -: TE)) = (`FD7THS_CP_R_QN_R, `FD7THS_CP_R_QN_F);
      if(!TI && E && D) (posedge CP => (QN +: TE)) = (`FD7THS_CP_R_QN_R, `FD7THS_CP_R_QN_F);
      if(!TI && !E && IQ) (posedge CP => (QN +: TE)) = (`FD7THS_CP_R_QN_R, `FD7THS_CP_R_QN_F);
      if(TE) (posedge CP => (QN -: TI)) = (`FD7THS_CP_R_QN_R, `FD7THS_CP_R_QN_F);
      if(!IQ && !TE && D) (posedge CP => (QN -: E)) = (`FD7THS_CP_R_QN_R, `FD7THS_CP_R_QN_F);
      if(!D && !TE && IQ) (posedge CP => (QN +: E)) = (`FD7THS_CP_R_QN_R, `FD7THS_CP_R_QN_F);
      if(!TE && E) (posedge CP => (QN -: D)) = (`FD7THS_CP_R_QN_R, `FD7THS_CP_R_QN_F);

      if(!IQ && !E && TI) (posedge CP => (SO +: TE)) = (`FD7THS_CP_R_SO_R, `FD7THS_CP_R_SO_F);
      if(!D && E && TI) (posedge CP => (SO +: TE)) = (`FD7THS_CP_R_SO_R, `FD7THS_CP_R_SO_F);
      if(!TI && E && D) (posedge CP => (SO -: TE)) = (`FD7THS_CP_R_SO_R, `FD7THS_CP_R_SO_F);
      if(!TI && !E && IQ) (posedge CP => (SO -: TE)) = (`FD7THS_CP_R_SO_R, `FD7THS_CP_R_SO_F);
      if(TE) (posedge CP => (SO +: TI)) = (`FD7THS_CP_R_SO_R, `FD7THS_CP_R_SO_F);
      if(!IQ && !TE && D) (posedge CP => (SO +: E)) = (`FD7THS_CP_R_SO_R, `FD7THS_CP_R_SO_F);
      if(!D && !TE && IQ) (posedge CP => (SO -: E)) = (`FD7THS_CP_R_SO_R, `FD7THS_CP_R_SO_F);
      if(!TE && E) (posedge CP => (SO +: D)) = (`FD7THS_CP_R_SO_R, `FD7THS_CP_R_SO_F);
 
	$setuphold(posedge CP &&& AndTEXE_, posedge D, `FD7THS_D_CP_SETUP_posedge_posedge, `FD7THS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndTEXE_, negedge D, `FD7THS_D_CP_SETUP_negedge_posedge, `FD7THS_D_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TEX, posedge E, `FD7THS_E_CP_SETUP_posedge_posedge, `FD7THS_E_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TEX, negedge E, `FD7THS_E_CP_SETUP_negedge_posedge, `FD7THS_E_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FD7THS_TI_CP_SETUP_posedge_posedge, `FD7THS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FD7THS_TI_CP_SETUP_negedge_posedge, `FD7THS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& D_orTI, posedge TE, `FD7THS_TE_CP_SETUP_posedge_posedge, `FD7THS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& D_orTI, negedge TE, `FD7THS_TE_CP_SETUP_negedge_posedge, `FD7THS_TE_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD7THS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7THS_CP_PWH, 0, Notifier);
`else

      (posedge CP => (Q +: Mux21Mux21IQDE_TITE_)) = (`FD7THS_CP_R_Q_R, `FD7THS_CP_R_Q_F);
      (posedge CP => (QN -: Mux21Mux21IQDE_TITE_)) = (`FD7THS_CP_R_QN_R, `FD7THS_CP_R_QN_F);
 
      (posedge CP => (SO +: Mux21Mux21IQDE_TITE_)) = (`FD7THS_CP_R_SO_R, `FD7THS_CP_R_SO_F);
 
        $setuphold(posedge CP &&& AndTEXE_, posedge D, `FD7THS_D_CP_SETUP_posedge_posedge, `FD7THS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndTEXE_, negedge D, `FD7THS_D_CP_SETUP_negedge_posedge, `FD7THS_D_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge E, `FD7THS_E_CP_SETUP_posedge_posedge, `FD7THS_E_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge E, `FD7THS_E_CP_SETUP_negedge_posedge, `FD7THS_E_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD7THS_TI_CP_SETUP_posedge_posedge, `FD7THS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD7THS_TI_CP_SETUP_negedge_posedge, `FD7THS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& D_orTI, posedge TE, `FD7THS_TE_CP_SETUP_posedge_posedge, `FD7THS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& D_orTI, negedge TE, `FD7THS_TE_CP_SETUP_negedge_posedge, `FD7THS_TE_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD7THS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7THS_CP_PWH, 0, Notifier);
`endif
 
   endspecify
`endif
 
endmodule // FD7THS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:57 and Version :1.1 //
 
//  START 
// CELL FD7THSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD7THSP_CP_R_QN_F 0.1
`define FD7THSP_CP_R_QN_R 0.1
`define FD7THSP_CP_R_Q_R 0.1
`define FD7THSP_CP_R_Q_F 0.1
`define FD7THSP_CP_R_SO_R 0.1
`define FD7THSP_CP_R_SO_F 0.1
`define FD7THSP_CP_PWH 0.1
`define FD7THSP_CP_PWL 0.1
`define FD7THSP_TE_CP_SETUP_posedge_posedge 0.1
`define FD7THSP_TE_CP_SETUP_negedge_posedge 0.1
`define FD7THSP_TE_CP_HOLD_posedge_posedge 0.1
`define FD7THSP_TE_CP_HOLD_negedge_posedge 0.1
`define FD7THSP_TI_CP_SETUP_posedge_posedge 0.1
`define FD7THSP_TI_CP_SETUP_negedge_posedge 0.1
`define FD7THSP_TI_CP_HOLD_posedge_posedge 0.1
`define FD7THSP_TI_CP_HOLD_negedge_posedge 0.1
`define FD7THSP_E_CP_SETUP_posedge_posedge 0.1
`define FD7THSP_E_CP_SETUP_negedge_posedge 0.1
`define FD7THSP_E_CP_HOLD_posedge_posedge 0.1
`define FD7THSP_E_CP_HOLD_negedge_posedge 0.1
`define FD7THSP_D_CP_SETUP_posedge_posedge 0.1
`define FD7THSP_D_CP_SETUP_negedge_posedge 0.1
`define FD7THSP_D_CP_HOLD_posedge_posedge 0.1
`define FD7THSP_D_CP_HOLD_negedge_posedge 0.1
 
module FD7THSP (Q, QN, SO, D, E, CP, TI, TE);
 
   output Q;
   output QN;
   output SO;
   input CP;
   input TE;
   input TI;
   input E;
   input D;
 
 
   reg Notifier;
 
   U_MUX2  u0 (Mux21IQDE_, IQ, D, E);
   U_MUX2  u1 (Mux21Mux21IQDE_TITE_, Mux21IQDE_, TI, TE);
 
   U_FD_P_NOTI u2 (   // Verilog Seq UDP
     IQ, Mux21Mux21IQDE_TITE_, CP, Notifier);
 
   buf  u3 (Q, IQ);
   not  u4 (QN, IQ);
   buf  u5 (SO, IQ);
 
 
 
`ifdef functional
`else
   and  (DE_, D, E);
   and  (QE_, Q, E_);
    or  (DEor_, DE_, QE_);
   not  (E_, E);

   xor  (D_orTI, DEor_, TI);
   not  (TEX, TE);
   and  (AndTEXE_, TEX, E);
   specify
`ifdef verifault
 
      if(!IQ && !E && TI) (posedge CP => (Q +: TE)) = (`FD7THSP_CP_R_Q_R, `FD7THSP_CP_R_Q_F);
      if(!D && E && TI) (posedge CP => (Q +: TE)) = (`FD7THSP_CP_R_Q_R, `FD7THSP_CP_R_Q_F);
      if(!TI && E && D) (posedge CP => (Q -: TE)) = (`FD7THSP_CP_R_Q_R, `FD7THSP_CP_R_Q_F);
      if(!TI && !E && IQ) (posedge CP => (Q -: TE)) = (`FD7THSP_CP_R_Q_R, `FD7THSP_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD7THSP_CP_R_Q_R, `FD7THSP_CP_R_Q_F);
      if(!IQ && !TE && D) (posedge CP => (Q +: E)) = (`FD7THSP_CP_R_Q_R, `FD7THSP_CP_R_Q_F);
      if(!D && !TE && IQ) (posedge CP => (Q -: E)) = (`FD7THSP_CP_R_Q_R, `FD7THSP_CP_R_Q_F);
      if(!TE && E) (posedge CP => (Q +: D)) = (`FD7THSP_CP_R_Q_R, `FD7THSP_CP_R_Q_F);
      if(!IQ && !E && TI) (posedge CP => (QN -: TE)) = (`FD7THSP_CP_R_QN_R, `FD7THSP_CP_R_QN_F);
      if(!D && E && TI) (posedge CP => (QN -: TE)) = (`FD7THSP_CP_R_QN_R, `FD7THSP_CP_R_QN_F);
      if(!TI && E && D) (posedge CP => (QN +: TE)) = (`FD7THSP_CP_R_QN_R, `FD7THSP_CP_R_QN_F);
      if(!TI && !E && IQ) (posedge CP => (QN +: TE)) = (`FD7THSP_CP_R_QN_R, `FD7THSP_CP_R_QN_F);
      if(TE) (posedge CP => (QN -: TI)) = (`FD7THSP_CP_R_QN_R, `FD7THSP_CP_R_QN_F);
      if(!IQ && !TE && D) (posedge CP => (QN -: E)) = (`FD7THSP_CP_R_QN_R, `FD7THSP_CP_R_QN_F);
      if(!D && !TE && IQ) (posedge CP => (QN +: E)) = (`FD7THSP_CP_R_QN_R, `FD7THSP_CP_R_QN_F);
      if(!TE && E) (posedge CP => (QN -: D)) = (`FD7THSP_CP_R_QN_R, `FD7THSP_CP_R_QN_F);

      if(!IQ && !E && TI) (posedge CP => (SO +: TE)) = (`FD7THSP_CP_R_SO_R, `FD7THSP_CP_R_SO_F);
      if(!D && E && TI) (posedge CP => (SO +: TE)) = (`FD7THSP_CP_R_SO_R, `FD7THSP_CP_R_SO_F);
      if(!TI && E && D) (posedge CP => (SO -: TE)) = (`FD7THSP_CP_R_SO_R, `FD7THSP_CP_R_SO_F);
      if(!TI && !E && IQ) (posedge CP => (SO -: TE)) = (`FD7THSP_CP_R_SO_R, `FD7THSP_CP_R_SO_F);
      if(TE) (posedge CP => (SO +: TI)) = (`FD7THSP_CP_R_SO_R, `FD7THSP_CP_R_SO_F);
      if(!IQ && !TE && D) (posedge CP => (SO +: E)) = (`FD7THSP_CP_R_SO_R, `FD7THSP_CP_R_SO_F);
      if(!D && !TE && IQ) (posedge CP => (SO -: E)) = (`FD7THSP_CP_R_SO_R, `FD7THSP_CP_R_SO_F);
      if(!TE && E) (posedge CP => (SO +: D)) = (`FD7THSP_CP_R_SO_R, `FD7THSP_CP_R_SO_F);
 
	$setuphold(posedge CP &&& AndTEXE_, posedge D, `FD7THSP_D_CP_SETUP_posedge_posedge, `FD7THSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndTEXE_, negedge D, `FD7THSP_D_CP_SETUP_negedge_posedge, `FD7THSP_D_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TEX, posedge E, `FD7THSP_E_CP_SETUP_posedge_posedge, `FD7THSP_E_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TEX, negedge E, `FD7THSP_E_CP_SETUP_negedge_posedge, `FD7THSP_E_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FD7THSP_TI_CP_SETUP_posedge_posedge, `FD7THSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FD7THSP_TI_CP_SETUP_negedge_posedge, `FD7THSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& D_orTI, posedge TE, `FD7THSP_TE_CP_SETUP_posedge_posedge, `FD7THSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& D_orTI, negedge TE, `FD7THSP_TE_CP_SETUP_negedge_posedge, `FD7THSP_TE_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD7THSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7THSP_CP_PWH, 0, Notifier);
`else

      (posedge CP => (Q +: Mux21Mux21IQDE_TITE_)) = (`FD7THSP_CP_R_Q_R, `FD7THSP_CP_R_Q_F);
      (posedge CP => (QN -: Mux21Mux21IQDE_TITE_)) = (`FD7THSP_CP_R_QN_R, `FD7THSP_CP_R_QN_F);
 
      (posedge CP => (SO +: Mux21Mux21IQDE_TITE_)) = (`FD7THSP_CP_R_SO_R, `FD7THSP_CP_R_SO_F);
 
        $setuphold(posedge CP &&& AndTEXE_, posedge D, `FD7THSP_D_CP_SETUP_posedge_posedge, `FD7THSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndTEXE_, negedge D, `FD7THSP_D_CP_SETUP_negedge_posedge, `FD7THSP_D_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge E, `FD7THSP_E_CP_SETUP_posedge_posedge, `FD7THSP_E_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge E, `FD7THSP_E_CP_SETUP_negedge_posedge, `FD7THSP_E_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD7THSP_TI_CP_SETUP_posedge_posedge, `FD7THSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD7THSP_TI_CP_SETUP_negedge_posedge, `FD7THSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& D_orTI, posedge TE, `FD7THSP_TE_CP_SETUP_posedge_posedge, `FD7THSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& D_orTI, negedge TE, `FD7THSP_TE_CP_SETUP_negedge_posedge, `FD7THSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD7THSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7THSP_CP_PWH, 0, Notifier);
`endif
 
   endspecify
`endif
 
endmodule // FD7THSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:57 and Version :1.1 //
 
//  START 
// CELL FD7THSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD7THSX4_CP_R_QN_F 0.1
`define FD7THSX4_CP_R_QN_R 0.1
`define FD7THSX4_CP_R_Q_R 0.1
`define FD7THSX4_CP_R_Q_F 0.1
`define FD7THSX4_CP_R_SO_R 0.1
`define FD7THSX4_CP_R_SO_F 0.1
`define FD7THSX4_CP_PWH 0.1
`define FD7THSX4_CP_PWL 0.1
`define FD7THSX4_TE_CP_SETUP_posedge_posedge 0.1
`define FD7THSX4_TE_CP_SETUP_negedge_posedge 0.1
`define FD7THSX4_TE_CP_HOLD_posedge_posedge 0.1
`define FD7THSX4_TE_CP_HOLD_negedge_posedge 0.1
`define FD7THSX4_TI_CP_SETUP_posedge_posedge 0.1
`define FD7THSX4_TI_CP_SETUP_negedge_posedge 0.1
`define FD7THSX4_TI_CP_HOLD_posedge_posedge 0.1
`define FD7THSX4_TI_CP_HOLD_negedge_posedge 0.1
`define FD7THSX4_E_CP_SETUP_posedge_posedge 0.1
`define FD7THSX4_E_CP_SETUP_negedge_posedge 0.1
`define FD7THSX4_E_CP_HOLD_posedge_posedge 0.1
`define FD7THSX4_E_CP_HOLD_negedge_posedge 0.1
`define FD7THSX4_D_CP_SETUP_posedge_posedge 0.1
`define FD7THSX4_D_CP_SETUP_negedge_posedge 0.1
`define FD7THSX4_D_CP_HOLD_posedge_posedge 0.1
`define FD7THSX4_D_CP_HOLD_negedge_posedge 0.1
 
module FD7THSX4 (Q, QN, SO, D, E, CP, TI, TE);
 
   output Q;
   output QN;
   output SO;
   input CP;
   input TE;
   input TI;
   input E;
   input D;
 
 
   reg Notifier;
 
   U_MUX2  u0 (Mux21IQDE_, IQ, D, E);
   U_MUX2  u1 (Mux21Mux21IQDE_TITE_, Mux21IQDE_, TI, TE);
 
   U_FD_P_NOTI u2 (   // Verilog Seq UDP
     IQ, Mux21Mux21IQDE_TITE_, CP, Notifier);
 
   buf  u3 (Q, IQ);
   not  u4 (QN, IQ);
   buf  u5 (SO, IQ);
 
 
 
`ifdef functional
`else
   and  (DE_, D, E);
   and  (QE_, Q, E_);
    or  (DEor_, DE_, QE_);
   not  (E_, E);

   xor  (D_orTI, DEor_, TI);
   not  (TEX, TE);
   and  (AndTEXE_, TEX, E);
   specify
`ifdef verifault
 
      if(!IQ && !E && TI) (posedge CP => (Q +: TE)) = (`FD7THSX4_CP_R_Q_R, `FD7THSX4_CP_R_Q_F);
      if(!D && E && TI) (posedge CP => (Q +: TE)) = (`FD7THSX4_CP_R_Q_R, `FD7THSX4_CP_R_Q_F);
      if(!TI && E && D) (posedge CP => (Q -: TE)) = (`FD7THSX4_CP_R_Q_R, `FD7THSX4_CP_R_Q_F);
      if(!TI && !E && IQ) (posedge CP => (Q -: TE)) = (`FD7THSX4_CP_R_Q_R, `FD7THSX4_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD7THSX4_CP_R_Q_R, `FD7THSX4_CP_R_Q_F);
      if(!IQ && !TE && D) (posedge CP => (Q +: E)) = (`FD7THSX4_CP_R_Q_R, `FD7THSX4_CP_R_Q_F);
      if(!D && !TE && IQ) (posedge CP => (Q -: E)) = (`FD7THSX4_CP_R_Q_R, `FD7THSX4_CP_R_Q_F);
      if(!TE && E) (posedge CP => (Q +: D)) = (`FD7THSX4_CP_R_Q_R, `FD7THSX4_CP_R_Q_F);
      if(!IQ && !E && TI) (posedge CP => (QN -: TE)) = (`FD7THSX4_CP_R_QN_R, `FD7THSX4_CP_R_QN_F);
      if(!D && E && TI) (posedge CP => (QN -: TE)) = (`FD7THSX4_CP_R_QN_R, `FD7THSX4_CP_R_QN_F);
      if(!TI && E && D) (posedge CP => (QN +: TE)) = (`FD7THSX4_CP_R_QN_R, `FD7THSX4_CP_R_QN_F);
      if(!TI && !E && IQ) (posedge CP => (QN +: TE)) = (`FD7THSX4_CP_R_QN_R, `FD7THSX4_CP_R_QN_F);
      if(TE) (posedge CP => (QN -: TI)) = (`FD7THSX4_CP_R_QN_R, `FD7THSX4_CP_R_QN_F);
      if(!IQ && !TE && D) (posedge CP => (QN -: E)) = (`FD7THSX4_CP_R_QN_R, `FD7THSX4_CP_R_QN_F);
      if(!D && !TE && IQ) (posedge CP => (QN +: E)) = (`FD7THSX4_CP_R_QN_R, `FD7THSX4_CP_R_QN_F);
      if(!TE && E) (posedge CP => (QN -: D)) = (`FD7THSX4_CP_R_QN_R, `FD7THSX4_CP_R_QN_F);

      if(!IQ && !E && TI) (posedge CP => (SO +: TE)) = (`FD7THSX4_CP_R_SO_R, `FD7THSX4_CP_R_SO_F);
      if(!D && E && TI) (posedge CP => (SO +: TE)) = (`FD7THSX4_CP_R_SO_R, `FD7THSX4_CP_R_SO_F);
      if(!TI && E && D) (posedge CP => (SO -: TE)) = (`FD7THSX4_CP_R_SO_R, `FD7THSX4_CP_R_SO_F);
      if(!TI && !E && IQ) (posedge CP => (SO -: TE)) = (`FD7THSX4_CP_R_SO_R, `FD7THSX4_CP_R_SO_F);
      if(TE) (posedge CP => (SO +: TI)) = (`FD7THSX4_CP_R_SO_R, `FD7THSX4_CP_R_SO_F);
      if(!IQ && !TE && D) (posedge CP => (SO +: E)) = (`FD7THSX4_CP_R_SO_R, `FD7THSX4_CP_R_SO_F);
      if(!D && !TE && IQ) (posedge CP => (SO -: E)) = (`FD7THSX4_CP_R_SO_R, `FD7THSX4_CP_R_SO_F);
      if(!TE && E) (posedge CP => (SO +: D)) = (`FD7THSX4_CP_R_SO_R, `FD7THSX4_CP_R_SO_F);
 
	$setuphold(posedge CP &&& AndTEXE_, posedge D, `FD7THSX4_D_CP_SETUP_posedge_posedge, `FD7THSX4_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndTEXE_, negedge D, `FD7THSX4_D_CP_SETUP_negedge_posedge, `FD7THSX4_D_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TEX, posedge E, `FD7THSX4_E_CP_SETUP_posedge_posedge, `FD7THSX4_E_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TEX, negedge E, `FD7THSX4_E_CP_SETUP_negedge_posedge, `FD7THSX4_E_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FD7THSX4_TI_CP_SETUP_posedge_posedge, `FD7THSX4_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FD7THSX4_TI_CP_SETUP_negedge_posedge, `FD7THSX4_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& D_orTI, posedge TE, `FD7THSX4_TE_CP_SETUP_posedge_posedge, `FD7THSX4_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& D_orTI, negedge TE, `FD7THSX4_TE_CP_SETUP_negedge_posedge, `FD7THSX4_TE_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD7THSX4_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7THSX4_CP_PWH, 0, Notifier);
`else

      (posedge CP => (Q +: Mux21Mux21IQDE_TITE_)) = (`FD7THSX4_CP_R_Q_R, `FD7THSX4_CP_R_Q_F);
      (posedge CP => (QN -: Mux21Mux21IQDE_TITE_)) = (`FD7THSX4_CP_R_QN_R, `FD7THSX4_CP_R_QN_F);
 
      (posedge CP => (SO +: Mux21Mux21IQDE_TITE_)) = (`FD7THSX4_CP_R_SO_R, `FD7THSX4_CP_R_SO_F);
 
        $setuphold(posedge CP &&& AndTEXE_, posedge D, `FD7THSX4_D_CP_SETUP_posedge_posedge, `FD7THSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndTEXE_, negedge D, `FD7THSX4_D_CP_SETUP_negedge_posedge, `FD7THSX4_D_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge E, `FD7THSX4_E_CP_SETUP_posedge_posedge, `FD7THSX4_E_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge E, `FD7THSX4_E_CP_SETUP_negedge_posedge, `FD7THSX4_E_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD7THSX4_TI_CP_SETUP_posedge_posedge, `FD7THSX4_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD7THSX4_TI_CP_SETUP_negedge_posedge, `FD7THSX4_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& D_orTI, posedge TE, `FD7THSX4_TE_CP_SETUP_posedge_posedge, `FD7THSX4_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& D_orTI, negedge TE, `FD7THSX4_TE_CP_SETUP_negedge_posedge, `FD7THSX4_TE_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD7THSX4_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7THSX4_CP_PWH, 0, Notifier);
`endif
 
   endspecify
`endif
 
endmodule // FD7THSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:16:57 and Version :1.1 //
 
//  START 
// CELL FD7TQHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD7TQHS_CP_R_Q_R 0.1
`define FD7TQHS_CP_R_Q_F 0.1
`define FD7TQHS_CP_R_SO_R 0.1
`define FD7TQHS_CP_R_SO_F 0.1
`define FD7TQHS_CP_PWH 0.1
`define FD7TQHS_CP_PWL 0.1
`define FD7TQHS_TE_CP_SETUP_posedge_posedge 0.1
`define FD7TQHS_TE_CP_SETUP_negedge_posedge 0.1
`define FD7TQHS_TE_CP_HOLD_posedge_posedge 0.1
`define FD7TQHS_TE_CP_HOLD_negedge_posedge 0.1
`define FD7TQHS_TI_CP_SETUP_posedge_posedge 0.1
`define FD7TQHS_TI_CP_SETUP_negedge_posedge 0.1
`define FD7TQHS_TI_CP_HOLD_posedge_posedge 0.1
`define FD7TQHS_TI_CP_HOLD_negedge_posedge 0.1
`define FD7TQHS_E_CP_SETUP_posedge_posedge 0.1
`define FD7TQHS_E_CP_SETUP_negedge_posedge 0.1
`define FD7TQHS_E_CP_HOLD_posedge_posedge 0.1
`define FD7TQHS_E_CP_HOLD_negedge_posedge 0.1
`define FD7TQHS_D_CP_SETUP_posedge_posedge 0.1
`define FD7TQHS_D_CP_SETUP_negedge_posedge 0.1
`define FD7TQHS_D_CP_HOLD_posedge_posedge 0.1
`define FD7TQHS_D_CP_HOLD_negedge_posedge 0.1
 
module FD7TQHS (Q, SO, D, E, CP, TI, TE);
 
   output Q;
   output SO;
   input CP;
   input TE;
   input TI;
   input E;
   input D;
 
 
   reg Notifier;
 
   U_MUX2  u0 (Mux21IQDE_, IQ, D, E);
   U_MUX2  u1 (Mux21Mux21IQDE_TITE_, Mux21IQDE_, TI, TE);
 
   U_FD_P_NOTI u2 (   // Verilog Seq UDP
      IQ, Mux21Mux21IQDE_TITE_, CP, Notifier);
 
   buf  u3 (Q, IQ);
   buf  u4 (SO, IQ);
 
 
 
`ifdef functional
`else
   and  (DE_, D, E);
   and  (QE_, Q, E_);
    or  (DEor_, DE_, QE_);
   not  (E_, E);

   xor  (D_orTI, DEor_, TI);
   not  (TEX, TE);
   and  (AndTEXE_, TEX, E);
   specify
`ifdef verifault
 
      if(!IQ && !E && TI) (posedge CP => (Q +: TE)) = (`FD7TQHS_CP_R_Q_R, `FD7TQHS_CP_R_Q_F);
      if(!D && E && TI) (posedge CP => (Q +: TE)) = (`FD7TQHS_CP_R_Q_R, `FD7TQHS_CP_R_Q_F);
      if(!TI && E && D) (posedge CP => (Q -: TE)) = (`FD7TQHS_CP_R_Q_R, `FD7TQHS_CP_R_Q_F);
      if(!TI && !E && IQ) (posedge CP => (Q -: TE)) = (`FD7TQHS_CP_R_Q_R, `FD7TQHS_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD7TQHS_CP_R_Q_R, `FD7TQHS_CP_R_Q_F);
      if(!IQ && !TE && D) (posedge CP => (Q +: E)) = (`FD7TQHS_CP_R_Q_R, `FD7TQHS_CP_R_Q_F);
      if(!D && !TE && IQ) (posedge CP => (Q -: E)) = (`FD7TQHS_CP_R_Q_R, `FD7TQHS_CP_R_Q_F);
      if(!TE && E) (posedge CP => (Q +: D)) = (`FD7TQHS_CP_R_Q_R, `FD7TQHS_CP_R_Q_F);
 
      if(!IQ && !E && TI) (posedge CP => (SO +: TE)) = (`FD7TQHS_CP_R_SO_R, `FD7TQHS_CP_R_SO_F);
      if(!D && E && TI) (posedge CP => (SO +: TE)) = (`FD7TQHS_CP_R_SO_R, `FD7TQHS_CP_R_SO_F);
      if(!TI && E && D) (posedge CP => (SO -: TE)) = (`FD7TQHS_CP_R_SO_R, `FD7TQHS_CP_R_SO_F);
      if(!TI && !E && IQ) (posedge CP => (SO -: TE)) = (`FD7TQHS_CP_R_SO_R, `FD7TQHS_CP_R_SO_F);
      if(TE) (posedge CP => (SO +: TI)) = (`FD7TQHS_CP_R_SO_R, `FD7TQHS_CP_R_SO_F);
      if(!IQ && !TE && D) (posedge CP => (SO +: E)) = (`FD7TQHS_CP_R_SO_R, `FD7TQHS_CP_R_SO_F);
      if(!D && !TE && IQ) (posedge CP => (SO -: E)) = (`FD7TQHS_CP_R_SO_R, `FD7TQHS_CP_R_SO_F);
      if(!TE && E) (posedge CP => (SO +: D)) = (`FD7TQHS_CP_R_SO_R, `FD7TQHS_CP_R_SO_F);

	$setuphold(posedge CP &&& AndTEXE_, posedge D, `FD7TQHS_D_CP_SETUP_posedge_posedge, `FD7TQHS_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndTEXE_, negedge D, `FD7TQHS_D_CP_SETUP_negedge_posedge, `FD7TQHS_D_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TEX, posedge E, `FD7TQHS_E_CP_SETUP_posedge_posedge, `FD7TQHS_E_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TEX, negedge E, `FD7TQHS_E_CP_SETUP_negedge_posedge, `FD7TQHS_E_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FD7TQHS_TI_CP_SETUP_posedge_posedge, `FD7TQHS_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FD7TQHS_TI_CP_SETUP_negedge_posedge, `FD7TQHS_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& D_orTI, posedge TE, `FD7TQHS_TE_CP_SETUP_posedge_posedge, `FD7TQHS_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& D_orTI, negedge TE, `FD7TQHS_TE_CP_SETUP_negedge_posedge, `FD7TQHS_TE_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD7TQHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7TQHS_CP_PWH, 0, Notifier);
`else
      (posedge CP => (Q +: Mux21Mux21IQDE_TITE_)) = (`FD7TQHS_CP_R_Q_R, `FD7TQHS_CP_R_Q_F);
      (posedge CP => (SO +: Mux21Mux21IQDE_TITE_)) = (`FD7TQHS_CP_R_SO_R, `FD7TQHS_CP_R_SO_F);
 
        $setuphold(posedge CP &&& AndTEXE_, posedge D, `FD7TQHS_D_CP_SETUP_posedge_posedge, `FD7TQHS_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndTEXE_, negedge D, `FD7TQHS_D_CP_SETUP_negedge_posedge, `FD7TQHS_D_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge E, `FD7TQHS_E_CP_SETUP_posedge_posedge, `FD7TQHS_E_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge E, `FD7TQHS_E_CP_SETUP_negedge_posedge, `FD7TQHS_E_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD7TQHS_TI_CP_SETUP_posedge_posedge, `FD7TQHS_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD7TQHS_TI_CP_SETUP_negedge_posedge, `FD7TQHS_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& D_orTI, posedge TE, `FD7TQHS_TE_CP_SETUP_posedge_posedge, `FD7TQHS_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& D_orTI, negedge TE, `FD7TQHS_TE_CP_SETUP_negedge_posedge, `FD7TQHS_TE_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD7TQHS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7TQHS_CP_PWH, 0, Notifier);

`endif 
   endspecify
`endif
 
 
endmodule // FD7TQHS 
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:01 and Version :1.1 //
 
//  START 
// CELL FD7TQHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD7TQHSP_CP_R_Q_R 0.1
`define FD7TQHSP_CP_R_Q_F 0.1
`define FD7TQHSP_CP_R_SO_R 0.1
`define FD7TQHSP_CP_R_SO_F 0.1
`define FD7TQHSP_CP_PWH 0.1
`define FD7TQHSP_CP_PWL 0.1
`define FD7TQHSP_TE_CP_SETUP_posedge_posedge 0.1
`define FD7TQHSP_TE_CP_SETUP_negedge_posedge 0.1
`define FD7TQHSP_TE_CP_HOLD_posedge_posedge 0.1
`define FD7TQHSP_TE_CP_HOLD_negedge_posedge 0.1
`define FD7TQHSP_TI_CP_SETUP_posedge_posedge 0.1
`define FD7TQHSP_TI_CP_SETUP_negedge_posedge 0.1
`define FD7TQHSP_TI_CP_HOLD_posedge_posedge 0.1
`define FD7TQHSP_TI_CP_HOLD_negedge_posedge 0.1
`define FD7TQHSP_E_CP_SETUP_posedge_posedge 0.1
`define FD7TQHSP_E_CP_SETUP_negedge_posedge 0.1
`define FD7TQHSP_E_CP_HOLD_posedge_posedge 0.1
`define FD7TQHSP_E_CP_HOLD_negedge_posedge 0.1
`define FD7TQHSP_D_CP_SETUP_posedge_posedge 0.1
`define FD7TQHSP_D_CP_SETUP_negedge_posedge 0.1
`define FD7TQHSP_D_CP_HOLD_posedge_posedge 0.1
`define FD7TQHSP_D_CP_HOLD_negedge_posedge 0.1
 
module FD7TQHSP (Q, SO, D, E, CP, TI, TE);
 
   output Q;
   output SO;
   input CP;
   input TE;
   input TI;
   input E;
   input D;
 
 
   reg Notifier;
 
   U_MUX2  u0 (Mux21IQDE_, IQ, D, E);
   U_MUX2  u1 (Mux21Mux21IQDE_TITE_, Mux21IQDE_, TI, TE);
 
   U_FD_P_NOTI u2 (   // Verilog Seq UDP
      IQ, Mux21Mux21IQDE_TITE_, CP, Notifier);
 
   buf  u3 (Q, IQ);
   buf  u4 (SO, IQ);
 
 
 
`ifdef functional
`else
   and  (DE_, D, E);
   and  (QE_, Q, E_);
    or  (DEor_, DE_, QE_);
   not  (E_, E);

   xor  (D_orTI, DEor_, TI);
   not  (TEX, TE);
   and  (AndTEXE_, TEX, E);
   specify
`ifdef verifault
 
      if(!IQ && !E && TI) (posedge CP => (Q +: TE)) = (`FD7TQHSP_CP_R_Q_R, `FD7TQHSP_CP_R_Q_F);
      if(!D && E && TI) (posedge CP => (Q +: TE)) = (`FD7TQHSP_CP_R_Q_R, `FD7TQHSP_CP_R_Q_F);
      if(!TI && E && D) (posedge CP => (Q -: TE)) = (`FD7TQHSP_CP_R_Q_R, `FD7TQHSP_CP_R_Q_F);
      if(!TI && !E && IQ) (posedge CP => (Q -: TE)) = (`FD7TQHSP_CP_R_Q_R, `FD7TQHSP_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD7TQHSP_CP_R_Q_R, `FD7TQHSP_CP_R_Q_F);
      if(!IQ && !TE && D) (posedge CP => (Q +: E)) = (`FD7TQHSP_CP_R_Q_R, `FD7TQHSP_CP_R_Q_F);
      if(!D && !TE && IQ) (posedge CP => (Q -: E)) = (`FD7TQHSP_CP_R_Q_R, `FD7TQHSP_CP_R_Q_F);
      if(!TE && E) (posedge CP => (Q +: D)) = (`FD7TQHSP_CP_R_Q_R, `FD7TQHSP_CP_R_Q_F);
 
      if(!IQ && !E && TI) (posedge CP => (SO +: TE)) = (`FD7TQHSP_CP_R_SO_R, `FD7TQHSP_CP_R_SO_F);
      if(!D && E && TI) (posedge CP => (SO +: TE)) = (`FD7TQHSP_CP_R_SO_R, `FD7TQHSP_CP_R_SO_F);
      if(!TI && E && D) (posedge CP => (SO -: TE)) = (`FD7TQHSP_CP_R_SO_R, `FD7TQHSP_CP_R_SO_F);
      if(!TI && !E && IQ) (posedge CP => (SO -: TE)) = (`FD7TQHSP_CP_R_SO_R, `FD7TQHSP_CP_R_SO_F);
      if(TE) (posedge CP => (SO +: TI)) = (`FD7TQHSP_CP_R_SO_R, `FD7TQHSP_CP_R_SO_F);
      if(!IQ && !TE && D) (posedge CP => (SO +: E)) = (`FD7TQHSP_CP_R_SO_R, `FD7TQHSP_CP_R_SO_F);
      if(!D && !TE && IQ) (posedge CP => (SO -: E)) = (`FD7TQHSP_CP_R_SO_R, `FD7TQHSP_CP_R_SO_F);
      if(!TE && E) (posedge CP => (SO +: D)) = (`FD7TQHSP_CP_R_SO_R, `FD7TQHSP_CP_R_SO_F);

	$setuphold(posedge CP &&& AndTEXE_, posedge D, `FD7TQHSP_D_CP_SETUP_posedge_posedge, `FD7TQHSP_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndTEXE_, negedge D, `FD7TQHSP_D_CP_SETUP_negedge_posedge, `FD7TQHSP_D_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TEX, posedge E, `FD7TQHSP_E_CP_SETUP_posedge_posedge, `FD7TQHSP_E_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TEX, negedge E, `FD7TQHSP_E_CP_SETUP_negedge_posedge, `FD7TQHSP_E_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FD7TQHSP_TI_CP_SETUP_posedge_posedge, `FD7TQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FD7TQHSP_TI_CP_SETUP_negedge_posedge, `FD7TQHSP_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& D_orTI, posedge TE, `FD7TQHSP_TE_CP_SETUP_posedge_posedge, `FD7TQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& D_orTI, negedge TE, `FD7TQHSP_TE_CP_SETUP_negedge_posedge, `FD7TQHSP_TE_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD7TQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7TQHSP_CP_PWH, 0, Notifier);
`else
      (posedge CP => (Q +: Mux21Mux21IQDE_TITE_)) = (`FD7TQHSP_CP_R_Q_R, `FD7TQHSP_CP_R_Q_F);
      (posedge CP => (SO +: Mux21Mux21IQDE_TITE_)) = (`FD7TQHSP_CP_R_SO_R, `FD7TQHSP_CP_R_SO_F);
 
        $setuphold(posedge CP &&& AndTEXE_, posedge D, `FD7TQHSP_D_CP_SETUP_posedge_posedge, `FD7TQHSP_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndTEXE_, negedge D, `FD7TQHSP_D_CP_SETUP_negedge_posedge, `FD7TQHSP_D_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge E, `FD7TQHSP_E_CP_SETUP_posedge_posedge, `FD7TQHSP_E_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge E, `FD7TQHSP_E_CP_SETUP_negedge_posedge, `FD7TQHSP_E_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD7TQHSP_TI_CP_SETUP_posedge_posedge, `FD7TQHSP_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD7TQHSP_TI_CP_SETUP_negedge_posedge, `FD7TQHSP_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& D_orTI, posedge TE, `FD7TQHSP_TE_CP_SETUP_posedge_posedge, `FD7TQHSP_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& D_orTI, negedge TE, `FD7TQHSP_TE_CP_SETUP_negedge_posedge, `FD7TQHSP_TE_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD7TQHSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7TQHSP_CP_PWH, 0, Notifier);

`endif 
   endspecify
`endif
 
 
endmodule // FD7TQHSP 
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:01 and Version :1.1 //
 
//  START 
// CELL FD7TQHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FD7TQHSX4_CP_R_Q_R 0.1
`define FD7TQHSX4_CP_R_Q_F 0.1
`define FD7TQHSX4_CP_R_SO_R 0.1
`define FD7TQHSX4_CP_R_SO_F 0.1
`define FD7TQHSX4_CP_PWH 0.1
`define FD7TQHSX4_CP_PWL 0.1
`define FD7TQHSX4_TE_CP_SETUP_posedge_posedge 0.1
`define FD7TQHSX4_TE_CP_SETUP_negedge_posedge 0.1
`define FD7TQHSX4_TE_CP_HOLD_posedge_posedge 0.1
`define FD7TQHSX4_TE_CP_HOLD_negedge_posedge 0.1
`define FD7TQHSX4_TI_CP_SETUP_posedge_posedge 0.1
`define FD7TQHSX4_TI_CP_SETUP_negedge_posedge 0.1
`define FD7TQHSX4_TI_CP_HOLD_posedge_posedge 0.1
`define FD7TQHSX4_TI_CP_HOLD_negedge_posedge 0.1
`define FD7TQHSX4_E_CP_SETUP_posedge_posedge 0.1
`define FD7TQHSX4_E_CP_SETUP_negedge_posedge 0.1
`define FD7TQHSX4_E_CP_HOLD_posedge_posedge 0.1
`define FD7TQHSX4_E_CP_HOLD_negedge_posedge 0.1
`define FD7TQHSX4_D_CP_SETUP_posedge_posedge 0.1
`define FD7TQHSX4_D_CP_SETUP_negedge_posedge 0.1
`define FD7TQHSX4_D_CP_HOLD_posedge_posedge 0.1
`define FD7TQHSX4_D_CP_HOLD_negedge_posedge 0.1
 
module FD7TQHSX4 (Q, SO, D, E, CP, TI, TE);
 
   output Q;
   output SO;
   input CP;
   input TE;
   input TI;
   input E;
   input D;
 
 
   reg Notifier;
 
   U_MUX2  u0 (Mux21IQDE_, IQ, D, E);
   U_MUX2  u1 (Mux21Mux21IQDE_TITE_, Mux21IQDE_, TI, TE);
 
   U_FD_P_NOTI u2 (   // Verilog Seq UDP
      IQ, Mux21Mux21IQDE_TITE_, CP, Notifier);
 
   buf  u3 (Q, IQ);
   buf  u4 (SO, IQ);
 
 
 
`ifdef functional
`else
   and  (DE_, D, E);
   and  (QE_, Q, E_);
    or  (DEor_, DE_, QE_);
   not  (E_, E);

   xor  (D_orTI, DEor_, TI);
   not  (TEX, TE);
   and  (AndTEXE_, TEX, E);
   specify
`ifdef verifault
 
      if(!IQ && !E && TI) (posedge CP => (Q +: TE)) = (`FD7TQHSX4_CP_R_Q_R, `FD7TQHSX4_CP_R_Q_F);
      if(!D && E && TI) (posedge CP => (Q +: TE)) = (`FD7TQHSX4_CP_R_Q_R, `FD7TQHSX4_CP_R_Q_F);
      if(!TI && E && D) (posedge CP => (Q -: TE)) = (`FD7TQHSX4_CP_R_Q_R, `FD7TQHSX4_CP_R_Q_F);
      if(!TI && !E && IQ) (posedge CP => (Q -: TE)) = (`FD7TQHSX4_CP_R_Q_R, `FD7TQHSX4_CP_R_Q_F);
      if(TE) (posedge CP => (Q +: TI)) = (`FD7TQHSX4_CP_R_Q_R, `FD7TQHSX4_CP_R_Q_F);
      if(!IQ && !TE && D) (posedge CP => (Q +: E)) = (`FD7TQHSX4_CP_R_Q_R, `FD7TQHSX4_CP_R_Q_F);
      if(!D && !TE && IQ) (posedge CP => (Q -: E)) = (`FD7TQHSX4_CP_R_Q_R, `FD7TQHSX4_CP_R_Q_F);
      if(!TE && E) (posedge CP => (Q +: D)) = (`FD7TQHSX4_CP_R_Q_R, `FD7TQHSX4_CP_R_Q_F);
 
      if(!IQ && !E && TI) (posedge CP => (SO +: TE)) = (`FD7TQHSX4_CP_R_SO_R, `FD7TQHSX4_CP_R_SO_F);
      if(!D && E && TI) (posedge CP => (SO +: TE)) = (`FD7TQHSX4_CP_R_SO_R, `FD7TQHSX4_CP_R_SO_F);
      if(!TI && E && D) (posedge CP => (SO -: TE)) = (`FD7TQHSX4_CP_R_SO_R, `FD7TQHSX4_CP_R_SO_F);
      if(!TI && !E && IQ) (posedge CP => (SO -: TE)) = (`FD7TQHSX4_CP_R_SO_R, `FD7TQHSX4_CP_R_SO_F);
      if(TE) (posedge CP => (SO +: TI)) = (`FD7TQHSX4_CP_R_SO_R, `FD7TQHSX4_CP_R_SO_F);
      if(!IQ && !TE && D) (posedge CP => (SO +: E)) = (`FD7TQHSX4_CP_R_SO_R, `FD7TQHSX4_CP_R_SO_F);
      if(!D && !TE && IQ) (posedge CP => (SO -: E)) = (`FD7TQHSX4_CP_R_SO_R, `FD7TQHSX4_CP_R_SO_F);
      if(!TE && E) (posedge CP => (SO +: D)) = (`FD7TQHSX4_CP_R_SO_R, `FD7TQHSX4_CP_R_SO_F);

	$setuphold(posedge CP &&& AndTEXE_, posedge D, `FD7TQHSX4_D_CP_SETUP_posedge_posedge, `FD7TQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndTEXE_, negedge D, `FD7TQHSX4_D_CP_SETUP_negedge_posedge, `FD7TQHSX4_D_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TEX, posedge E, `FD7TQHSX4_E_CP_SETUP_posedge_posedge, `FD7TQHSX4_E_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TEX, negedge E, `FD7TQHSX4_E_CP_SETUP_negedge_posedge, `FD7TQHSX4_E_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& TE, posedge TI, `FD7TQHSX4_TI_CP_SETUP_posedge_posedge, `FD7TQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& TE, negedge TI, `FD7TQHSX4_TI_CP_SETUP_negedge_posedge, `FD7TQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& D_orTI, posedge TE, `FD7TQHSX4_TE_CP_SETUP_posedge_posedge, `FD7TQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& D_orTI, negedge TE, `FD7TQHSX4_TE_CP_SETUP_negedge_posedge, `FD7TQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FD7TQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7TQHSX4_CP_PWH, 0, Notifier);
`else
      (posedge CP => (Q +: Mux21Mux21IQDE_TITE_)) = (`FD7TQHSX4_CP_R_Q_R, `FD7TQHSX4_CP_R_Q_F);
      (posedge CP => (SO +: Mux21Mux21IQDE_TITE_)) = (`FD7TQHSX4_CP_R_SO_R, `FD7TQHSX4_CP_R_SO_F);
 
        $setuphold(posedge CP &&& AndTEXE_, posedge D, `FD7TQHSX4_D_CP_SETUP_posedge_posedge, `FD7TQHSX4_D_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndTEXE_, negedge D, `FD7TQHSX4_D_CP_SETUP_negedge_posedge, `FD7TQHSX4_D_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TEX, posedge E, `FD7TQHSX4_E_CP_SETUP_posedge_posedge, `FD7TQHSX4_E_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TEX, negedge E, `FD7TQHSX4_E_CP_SETUP_negedge_posedge, `FD7TQHSX4_E_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& TE, posedge TI, `FD7TQHSX4_TI_CP_SETUP_posedge_posedge, `FD7TQHSX4_TI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& TE, negedge TI, `FD7TQHSX4_TI_CP_SETUP_negedge_posedge, `FD7TQHSX4_TI_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& D_orTI, posedge TE, `FD7TQHSX4_TE_CP_SETUP_posedge_posedge, `FD7TQHSX4_TE_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& D_orTI, negedge TE, `FD7TQHSX4_TE_CP_SETUP_negedge_posedge, `FD7TQHSX4_TE_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FD7TQHSX4_CP_PWL, 0, Notifier);
      $width(posedge CP, `FD7TQHSX4_CP_PWH, 0, Notifier);

`endif 
   endspecify
`endif
 
 
endmodule // FD7TQHSX4 
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:01 and Version :1.1 //
 
//  START 
// CELL FJK1HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FJK1HS_CP_R_QN_R 0.1
`define FJK1HS_CP_R_QN_F 0.1
`define FJK1HS_CP_R_Q_F 0.1
`define FJK1HS_CP_R_Q_R 0.1
`define FJK1HS_CP_PWH 0.1
`define FJK1HS_CP_PWL 0.1
`define FJK1HS_J_CP_SETUP_posedge_posedge 0.1
`define FJK1HS_J_CP_SETUP_negedge_posedge 0.1
`define FJK1HS_J_CP_HOLD_posedge_posedge 0.1
`define FJK1HS_J_CP_HOLD_negedge_posedge 0.1
`define FJK1HS_K_CP_SETUP_posedge_posedge 0.1
`define FJK1HS_K_CP_SETUP_negedge_posedge 0.1
`define FJK1HS_K_CP_HOLD_posedge_posedge 0.1
`define FJK1HS_K_CP_HOLD_negedge_posedge 0.1

module FJK1HS (Q, QN, J, K, CP);

   output Q;
   output QN;
   input J;
   input K;
   input CP;


   reg Notifier;

   not  u0 (KX, K);
   U_MUX2  u1 (Mux21JKXIQ_, J, KX, IQ);

   U_FD_P_NOTI u2 (   // Verilog Seq UDP
      IQ, Mux21JKXIQ_, CP, Notifier);

   buf  u3 (Q, IQ);
   not  u4 (QN, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(!IQ) (posedge CP => (Q +: J)) = (`FJK1HS_CP_R_Q_R, `FJK1HS_CP_R_Q_F);
      if(IQ) (posedge CP => (Q -: K)) = (`FJK1HS_CP_R_Q_R, `FJK1HS_CP_R_Q_F);
      if(!IQ) (posedge CP => (QN -: J)) = (`FJK1HS_CP_R_QN_R, `FJK1HS_CP_R_QN_F);
      if(IQ) (posedge CP => (QN +: K)) = (`FJK1HS_CP_R_QN_R, `FJK1HS_CP_R_QN_F);

	$setuphold(posedge CP, posedge K, `FJK1HS_K_CP_SETUP_posedge_posedge, `FJK1HS_K_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP, negedge K, `FJK1HS_K_CP_SETUP_negedge_posedge, `FJK1HS_K_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP, posedge J, `FJK1HS_J_CP_SETUP_posedge_posedge, `FJK1HS_J_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP, negedge J, `FJK1HS_J_CP_SETUP_negedge_posedge, `FJK1HS_J_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FJK1HS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FJK1HS_CP_PWH, 0, Notifier);
`else

      (posedge CP => (Q +: Mux21JKXIQ_)) = (`FJK1HS_CP_R_Q_R, `FJK1HS_CP_R_Q_F);
      (posedge CP => (QN -: Mux21JKXIQ_)) = (`FJK1HS_CP_R_QN_R, `FJK1HS_CP_R_QN_F);
 
        $setuphold(posedge CP, posedge K, `FJK1HS_K_CP_SETUP_posedge_posedge, `FJK1HS_K_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP, negedge K, `FJK1HS_K_CP_SETUP_negedge_posedge, `FJK1HS_K_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP, posedge J, `FJK1HS_J_CP_SETUP_posedge_posedge, `FJK1HS_J_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP, negedge J, `FJK1HS_J_CP_SETUP_negedge_posedge, `FJK1HS_J_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FJK1HS_CP_PWL, 0, Notifier);
      $width(posedge CP, `FJK1HS_CP_PWH, 0, Notifier);
`endif
   endspecify
`endif


endmodule // FJK1HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:01 and Version :1.1 //
 
//  START 
// CELL FJK1HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FJK1HSP_CP_R_QN_R 0.1
`define FJK1HSP_CP_R_QN_F 0.1
`define FJK1HSP_CP_R_Q_F 0.1
`define FJK1HSP_CP_R_Q_R 0.1
`define FJK1HSP_CP_PWH 0.1
`define FJK1HSP_CP_PWL 0.1
`define FJK1HSP_J_CP_SETUP_posedge_posedge 0.1
`define FJK1HSP_J_CP_SETUP_negedge_posedge 0.1
`define FJK1HSP_J_CP_HOLD_posedge_posedge 0.1
`define FJK1HSP_J_CP_HOLD_negedge_posedge 0.1
`define FJK1HSP_K_CP_SETUP_posedge_posedge 0.1
`define FJK1HSP_K_CP_SETUP_negedge_posedge 0.1
`define FJK1HSP_K_CP_HOLD_posedge_posedge 0.1
`define FJK1HSP_K_CP_HOLD_negedge_posedge 0.1

module FJK1HSP (Q, QN, J, K, CP);

   output Q;
   output QN;
   input J;
   input K;
   input CP;


   reg Notifier;

   not  u0 (KX, K);
   U_MUX2  u1 (Mux21JKXIQ_, J, KX, IQ);

   U_FD_P_NOTI u2 (   // Verilog Seq UDP
      IQ, Mux21JKXIQ_, CP, Notifier);

   buf  u3 (Q, IQ);
   not  u4 (QN, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(!IQ) (posedge CP => (Q +: J)) = (`FJK1HSP_CP_R_Q_R, `FJK1HSP_CP_R_Q_F);
      if(IQ) (posedge CP => (Q -: K)) = (`FJK1HSP_CP_R_Q_R, `FJK1HSP_CP_R_Q_F);
      if(!IQ) (posedge CP => (QN -: J)) = (`FJK1HSP_CP_R_QN_R, `FJK1HSP_CP_R_QN_F);
      if(IQ) (posedge CP => (QN +: K)) = (`FJK1HSP_CP_R_QN_R, `FJK1HSP_CP_R_QN_F);

	$setuphold(posedge CP, posedge K, `FJK1HSP_K_CP_SETUP_posedge_posedge, `FJK1HSP_K_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP, negedge K, `FJK1HSP_K_CP_SETUP_negedge_posedge, `FJK1HSP_K_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP, posedge J, `FJK1HSP_J_CP_SETUP_posedge_posedge, `FJK1HSP_J_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP, negedge J, `FJK1HSP_J_CP_SETUP_negedge_posedge, `FJK1HSP_J_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FJK1HSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FJK1HSP_CP_PWH, 0, Notifier);
`else

      (posedge CP => (Q +: Mux21JKXIQ_)) = (`FJK1HSP_CP_R_Q_R, `FJK1HSP_CP_R_Q_F);
      (posedge CP => (QN -: Mux21JKXIQ_)) = (`FJK1HSP_CP_R_QN_R, `FJK1HSP_CP_R_QN_F);
 
        $setuphold(posedge CP, posedge K, `FJK1HSP_K_CP_SETUP_posedge_posedge, `FJK1HSP_K_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP, negedge K, `FJK1HSP_K_CP_SETUP_negedge_posedge, `FJK1HSP_K_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP, posedge J, `FJK1HSP_J_CP_SETUP_posedge_posedge, `FJK1HSP_J_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP, negedge J, `FJK1HSP_J_CP_SETUP_negedge_posedge, `FJK1HSP_J_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FJK1HSP_CP_PWL, 0, Notifier);
      $width(posedge CP, `FJK1HSP_CP_PWH, 0, Notifier);
`endif
   endspecify
`endif


endmodule // FJK1HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:01 and Version :1.1 //
 
//  START 
// CELL FJK2HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FJK2HS_CD_F_QN_R 0.1
`define FJK2HS_CP_R_QN_R 0.1
`define FJK2HS_CP_R_QN_F 0.1
`define FJK2HS_CD_F_Q_F 0.1
`define FJK2HS_CP_R_Q_F 0.1
`define FJK2HS_CP_R_Q_R 0.1
`define FJK2HS_CD_CP_REM_posedge_posedge 0.1
`define FJK2HS_CD_CP_REC_posedge_posedge 0.1
`define FJK2HS_CD_PWL 0.1
`define FJK2HS_CP_PWH 0.1
`define FJK2HS_CP_PWL 0.1
`define FJK2HS_J_CP_SETUP_posedge_posedge 0.1
`define FJK2HS_J_CP_SETUP_negedge_posedge 0.1
`define FJK2HS_J_CP_HOLD_posedge_posedge 0.1
`define FJK2HS_J_CP_HOLD_negedge_posedge 0.1
`define FJK2HS_K_CP_SETUP_posedge_posedge 0.1
`define FJK2HS_K_CP_SETUP_negedge_posedge 0.1
`define FJK2HS_K_CP_HOLD_posedge_posedge 0.1
`define FJK2HS_K_CP_HOLD_negedge_posedge 0.1

module FJK2HS (Q, QN, J, K, CP, CD);

   output Q;
   output QN;
   input J;
   input K;
   input CP;
   input CD;


   reg Notifier;

   not  u0 (KX, K);
   U_MUX2  u1 (Mux21JKXIQ_, J, KX, IQ);

   U_FD_P_RN_NOTI u2 ( IQ, Mux21JKXIQ_, CP, CD, Notifier);

   buf  u3 (Q, IQ);
   not  u4 (QN, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(!IQ) (posedge CP => (Q +: J)) = (`FJK2HS_CP_R_Q_R, `FJK2HS_CP_R_Q_F);
      if(IQ) (posedge CP => (Q -: K)) = (`FJK2HS_CP_R_Q_R, `FJK2HS_CP_R_Q_F);
      if(!IQ) (posedge CP => (QN -: J)) = (`FJK2HS_CP_R_QN_R, `FJK2HS_CP_R_QN_F);
      if(IQ) (posedge CP => (QN +: K)) = (`FJK2HS_CP_R_QN_R, `FJK2HS_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FJK2HS_CD_F_Q_F,`FJK2HS_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FJK2HS_CD_F_QN_R,`FJK2HS_CD_F_QN_R);

	$setuphold(posedge CP &&& CD, posedge K, `FJK2HS_K_CP_SETUP_posedge_posedge, `FJK2HS_K_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge K, `FJK2HS_K_CP_SETUP_negedge_posedge, `FJK2HS_K_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& CD, posedge J, `FJK2HS_J_CP_SETUP_posedge_posedge, `FJK2HS_J_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge J, `FJK2HS_J_CP_SETUP_negedge_posedge, `FJK2HS_J_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FJK2HS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FJK2HS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FJK2HS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& J, `FJK2HS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& J, posedge CD, `FJK2HS_CD_CP_REM_posedge_posedge, Notifier);

`else

      (posedge CP => (Q +: Mux21JKXIQ_)) = (`FJK2HS_CP_R_Q_R, `FJK2HS_CP_R_Q_F);
      (posedge CP => (QN -: Mux21JKXIQ_)) = (`FJK2HS_CP_R_QN_R, `FJK2HS_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FJK2HS_CD_F_Q_F,`FJK2HS_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FJK2HS_CD_F_QN_R,`FJK2HS_CD_F_QN_R);
 
        $setuphold(posedge CP &&& CD, posedge K, `FJK2HS_K_CP_SETUP_posedge_posedge, `FJK2HS_K_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge K, `FJK2HS_K_CP_SETUP_negedge_posedge, `FJK2HS_K_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& CD, posedge J, `FJK2HS_J_CP_SETUP_posedge_posedge, `FJK2HS_J_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge J, `FJK2HS_J_CP_SETUP_negedge_posedge, `FJK2HS_J_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FJK2HS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FJK2HS_CP_PWH, 0, Notifier);
      $width(negedge CD, `FJK2HS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& J, `FJK2HS_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& J, posedge CD, `FJK2HS_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FJK2HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:08 and Version :1.1 //
 
//  START 
// CELL FJK2HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FJK2HSP_CD_F_QN_R 0.1
`define FJK2HSP_CP_R_QN_R 0.1
`define FJK2HSP_CP_R_QN_F 0.1
`define FJK2HSP_CD_F_Q_F 0.1
`define FJK2HSP_CP_R_Q_F 0.1
`define FJK2HSP_CP_R_Q_R 0.1
`define FJK2HSP_CD_CP_REM_posedge_posedge 0.1
`define FJK2HSP_CD_CP_REC_posedge_posedge 0.1
`define FJK2HSP_CD_PWL 0.1
`define FJK2HSP_CP_PWH 0.1
`define FJK2HSP_CP_PWL 0.1
`define FJK2HSP_J_CP_SETUP_posedge_posedge 0.1
`define FJK2HSP_J_CP_SETUP_negedge_posedge 0.1
`define FJK2HSP_J_CP_HOLD_posedge_posedge 0.1
`define FJK2HSP_J_CP_HOLD_negedge_posedge 0.1
`define FJK2HSP_K_CP_SETUP_posedge_posedge 0.1
`define FJK2HSP_K_CP_SETUP_negedge_posedge 0.1
`define FJK2HSP_K_CP_HOLD_posedge_posedge 0.1
`define FJK2HSP_K_CP_HOLD_negedge_posedge 0.1

module FJK2HSP (Q, QN, J, K, CP, CD);

   output Q;
   output QN;
   input J;
   input K;
   input CP;
   input CD;


   reg Notifier;

   not  u0 (KX, K);
   U_MUX2  u1 (Mux21JKXIQ_, J, KX, IQ);

   U_FD_P_RN_NOTI u2 ( IQ, Mux21JKXIQ_, CP, CD, Notifier);

   buf  u3 (Q, IQ);
   not  u4 (QN, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(!IQ) (posedge CP => (Q +: J)) = (`FJK2HSP_CP_R_Q_R, `FJK2HSP_CP_R_Q_F);
      if(IQ) (posedge CP => (Q -: K)) = (`FJK2HSP_CP_R_Q_R, `FJK2HSP_CP_R_Q_F);
      if(!IQ) (posedge CP => (QN -: J)) = (`FJK2HSP_CP_R_QN_R, `FJK2HSP_CP_R_QN_F);
      if(IQ) (posedge CP => (QN +: K)) = (`FJK2HSP_CP_R_QN_R, `FJK2HSP_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FJK2HSP_CD_F_Q_F,`FJK2HSP_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FJK2HSP_CD_F_QN_R,`FJK2HSP_CD_F_QN_R);

	$setuphold(posedge CP &&& CD, posedge K, `FJK2HSP_K_CP_SETUP_posedge_posedge, `FJK2HSP_K_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge K, `FJK2HSP_K_CP_SETUP_negedge_posedge, `FJK2HSP_K_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& CD, posedge J, `FJK2HSP_J_CP_SETUP_posedge_posedge, `FJK2HSP_J_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge J, `FJK2HSP_J_CP_SETUP_negedge_posedge, `FJK2HSP_J_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FJK2HSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FJK2HSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `FJK2HSP_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP &&& J, `FJK2HSP_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& J, posedge CD, `FJK2HSP_CD_CP_REM_posedge_posedge, Notifier);

`else

      (posedge CP => (Q +: Mux21JKXIQ_)) = (`FJK2HSP_CP_R_Q_R, `FJK2HSP_CP_R_Q_F);
      (posedge CP => (QN -: Mux21JKXIQ_)) = (`FJK2HSP_CP_R_QN_R, `FJK2HSP_CP_R_QN_F);
      (negedge CD => (Q +: 1'b0)) = (`FJK2HSP_CD_F_Q_F,`FJK2HSP_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`FJK2HSP_CD_F_QN_R,`FJK2HSP_CD_F_QN_R);
 
        $setuphold(posedge CP &&& CD, posedge K, `FJK2HSP_K_CP_SETUP_posedge_posedge, `FJK2HSP_K_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge K, `FJK2HSP_K_CP_SETUP_negedge_posedge, `FJK2HSP_K_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& CD, posedge J, `FJK2HSP_J_CP_SETUP_posedge_posedge, `FJK2HSP_J_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge J, `FJK2HSP_J_CP_SETUP_negedge_posedge, `FJK2HSP_J_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FJK2HSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `FJK2HSP_CP_PWH, 0, Notifier);
      $width(negedge CD, `FJK2HSP_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP &&& J, `FJK2HSP_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& J, posedge CD, `FJK2HSP_CD_CP_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FJK2HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:08 and Version :1.1 //
 
//  START 
// CELL FJK3HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FJK3HS_SD_F_QN_F 0.1
`define FJK3HS_CD_F_QN_R 0.1
`define FJK3HS_CD_R_QN_F 0.1
`define FJK3HS_CP_R_QN_R 0.1
`define FJK3HS_CP_R_QN_F 0.1
`define FJK3HS_SD_F_Q_R 0.1
`define FJK3HS_CD_F_Q_F 0.1
`define FJK3HS_CD_R_Q_R 0.1
`define FJK3HS_CP_R_Q_F 0.1
`define FJK3HS_CP_R_Q_R 0.1
`define FJK3HS_CD_SD_REM_posedge_posedge 0.1
`define FJK3HS_CD_SD_REC_posedge_posedge 0.1
`define FJK3HS_CD_CP_REM_posedge_posedge 0.1
`define FJK3HS_SD_CP_REM_posedge_posedge 0.1
`define FJK3HS_CD_CP_REC_posedge_posedge 0.1
`define FJK3HS_SD_CP_REC_posedge_posedge 0.1
`define FJK3HS_CD_PWL 0.1
`define FJK3HS_SD_PWL 0.1
`define FJK3HS_CP_PWH 0.1
`define FJK3HS_CP_PWL 0.1
`define FJK3HS_J_CP_SETUP_posedge_posedge 0.1
`define FJK3HS_J_CP_SETUP_negedge_posedge 0.1
`define FJK3HS_J_CP_HOLD_posedge_posedge 0.1
`define FJK3HS_J_CP_HOLD_negedge_posedge 0.1
`define FJK3HS_K_CP_SETUP_posedge_posedge 0.1
`define FJK3HS_K_CP_SETUP_negedge_posedge 0.1
`define FJK3HS_K_CP_HOLD_posedge_posedge 0.1
`define FJK3HS_K_CP_HOLD_negedge_posedge 0.1

module FJK3HS (Q, QN, J, K, CP, CD, SD);

   output Q;
   output QN;
   input J;
   input K;
   input CP;
   input CD;
   input SD;


   reg Notifier;

   not  u0 (KX, K);
   U_MUX2  u1 (Mux21JKXIQ_, J, KX, IQ);

   U_FD_P_RN_SN_NOTI u2 (   // Verilog Seq UDP
      IQ, Mux21JKXIQ_, CP, CD, SD, Notifier);

   buf  u3 (Q, IQ);
   not  u4 (QN, IQ);



`ifdef functional
`else
   and  (AndCDSD_, CD, SD);
   and  (AndSDJ, SD, J);
   and  (AndCDK, CD, K);

   specify
`ifdef verifault

      if(!IQ && CD && SD) (posedge CP => (Q +: J)) = (`FJK3HS_CP_R_Q_R, `FJK3HS_CP_R_Q_F);
      if(IQ && CD && SD) (posedge CP => (Q -: K)) = (`FJK3HS_CP_R_Q_R, `FJK3HS_CP_R_Q_F);
      if(!IQ && CD && SD) (posedge CP => (QN -: J)) = (`FJK3HS_CP_R_QN_R, `FJK3HS_CP_R_QN_F);
      if(IQ && CD && SD) (posedge CP => (QN +: K)) = (`FJK3HS_CP_R_QN_R, `FJK3HS_CP_R_QN_F);
      if(!SD) (posedge CD => (Q +: 1'b1)) = (`FJK3HS_CD_R_Q_R,`FJK3HS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FJK3HS_CD_R_Q_R,`FJK3HS_CD_F_Q_F);
      if(CD) (negedge SD => (Q +: 1'b1)) = (`FJK3HS_SD_F_Q_R,`FJK3HS_SD_F_Q_R);
      if(!SD) (posedge CD => (QN +: 1'b0)) = (`FJK3HS_CD_F_QN_R,`FJK3HS_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`FJK3HS_CD_F_QN_R,`FJK3HS_CD_R_QN_F);
      if(CD) (negedge SD => (QN +: 1'b0)) = (`FJK3HS_SD_F_QN_F,`FJK3HS_SD_F_QN_F);

	$setuphold(posedge CP &&& AndCDSD_, posedge K, `FJK3HS_K_CP_SETUP_posedge_posedge, `FJK3HS_K_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSD_, negedge K, `FJK3HS_K_CP_SETUP_negedge_posedge, `FJK3HS_K_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDSD_, posedge J, `FJK3HS_J_CP_SETUP_posedge_posedge, `FJK3HS_J_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSD_, negedge J, `FJK3HS_J_CP_SETUP_negedge_posedge, `FJK3HS_J_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FJK3HS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FJK3HS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FJK3HS_SD_PWL, 0, Notifier);
      $width(negedge CD, `FJK3HS_CD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& AndCDK, `FJK3HS_SD_CP_REC_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge CP &&& AndSDJ, `FJK3HS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndCDK, posedge SD, `FJK3HS_SD_CP_REM_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndSDJ, posedge CD, `FJK3HS_CD_CP_REM_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge SD, `FJK3HS_CD_SD_REC_posedge_posedge, Notifier);

	$hold(posedge SD, posedge CD, `FJK3HS_CD_SD_REM_posedge_posedge, Notifier);

`else

      (posedge CP => (Q +: Mux21JKXIQ_)) = (`FJK3HS_CP_R_Q_R, `FJK3HS_CP_R_Q_F);
      (posedge CP => (QN -: Mux21JKXIQ_)) = (`FJK3HS_CP_R_QN_R, `FJK3HS_CP_R_QN_F);
      (posedge CD => (Q +: 1'b1)) = (`FJK3HS_CD_R_Q_R,`FJK3HS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FJK3HS_CD_R_Q_R,`FJK3HS_CD_F_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FJK3HS_SD_F_Q_R,`FJK3HS_SD_F_Q_R);
      (posedge CD => (QN +: 1'b0)) = (`FJK3HS_CD_F_QN_R,`FJK3HS_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`FJK3HS_CD_F_QN_R,`FJK3HS_CD_R_QN_F);
      (negedge SD => (QN +: 1'b0)) = (`FJK3HS_SD_F_QN_F,`FJK3HS_SD_F_QN_F);
 
        $setuphold(posedge CP &&& AndCDSD_, posedge K, `FJK3HS_K_CP_SETUP_posedge_posedge, `FJK3HS_K_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSD_, negedge K, `FJK3HS_K_CP_SETUP_negedge_posedge, `FJK3HS_K_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDSD_, posedge J, `FJK3HS_J_CP_SETUP_posedge_posedge, `FJK3HS_J_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSD_, negedge J, `FJK3HS_J_CP_SETUP_negedge_posedge, `FJK3HS_J_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FJK3HS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FJK3HS_CP_PWH, 0, Notifier);
      $width(negedge SD, `FJK3HS_SD_PWL, 0, Notifier);
      $width(negedge CD, `FJK3HS_CD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& AndCDK, `FJK3HS_SD_CP_REC_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge CP &&& AndSDJ, `FJK3HS_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndCDK, posedge SD, `FJK3HS_SD_CP_REM_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndSDJ, posedge CD, `FJK3HS_CD_CP_REM_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge SD, `FJK3HS_CD_SD_REC_posedge_posedge, Notifier);
 
        $hold(posedge SD, posedge CD, `FJK3HS_CD_SD_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FJK3HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:15 and Version :1.1 //
 
//  START 
// CELL FJK3HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define FJK3HSP_SD_F_QN_F 0.1
`define FJK3HSP_CD_F_QN_R 0.1
`define FJK3HSP_CD_R_QN_F 0.1
`define FJK3HSP_CP_R_QN_R 0.1
`define FJK3HSP_CP_R_QN_F 0.1
`define FJK3HSP_SD_F_Q_R 0.1
`define FJK3HSP_CD_F_Q_F 0.1
`define FJK3HSP_CD_R_Q_R 0.1
`define FJK3HSP_CP_R_Q_F 0.1
`define FJK3HSP_CP_R_Q_R 0.1
`define FJK3HSP_CD_SD_REM_posedge_posedge 0.1
`define FJK3HSP_CD_SD_REC_posedge_posedge 0.1
`define FJK3HSP_CD_CP_REM_posedge_posedge 0.1
`define FJK3HSP_SD_CP_REM_posedge_posedge 0.1
`define FJK3HSP_CD_CP_REC_posedge_posedge 0.1
`define FJK3HSP_SD_CP_REC_posedge_posedge 0.1
`define FJK3HSP_CD_PWL 0.1
`define FJK3HSP_SD_PWL 0.1
`define FJK3HSP_CP_PWH 0.1
`define FJK3HSP_CP_PWL 0.1
`define FJK3HSP_J_CP_SETUP_posedge_posedge 0.1
`define FJK3HSP_J_CP_SETUP_negedge_posedge 0.1
`define FJK3HSP_J_CP_HOLD_posedge_posedge 0.1
`define FJK3HSP_J_CP_HOLD_negedge_posedge 0.1
`define FJK3HSP_K_CP_SETUP_posedge_posedge 0.1
`define FJK3HSP_K_CP_SETUP_negedge_posedge 0.1
`define FJK3HSP_K_CP_HOLD_posedge_posedge 0.1
`define FJK3HSP_K_CP_HOLD_negedge_posedge 0.1

module FJK3HSP (Q, QN, J, K, CP, CD, SD);

   output Q;
   output QN;
   input J;
   input K;
   input CP;
   input CD;
   input SD;


   reg Notifier;

   not  u0 (KX, K);
   U_MUX2  u1 (Mux21JKXIQ_, J, KX, IQ);

   U_FD_P_RN_SN_NOTI u2 (   // Verilog Seq UDP
      IQ, Mux21JKXIQ_, CP, CD, SD, Notifier);

   buf  u3 (Q, IQ);
   not  u4 (QN, IQ);



`ifdef functional
`else
   and  (AndCDSD_, CD, SD);
   and  (AndSDJ, SD, J);
   and  (AndCDK, CD, K);

   specify
`ifdef verifault

      if(!IQ && CD && SD) (posedge CP => (Q +: J)) = (`FJK3HSP_CP_R_Q_R, `FJK3HSP_CP_R_Q_F);
      if(IQ && CD && SD) (posedge CP => (Q -: K)) = (`FJK3HSP_CP_R_Q_R, `FJK3HSP_CP_R_Q_F);
      if(!IQ && CD && SD) (posedge CP => (QN -: J)) = (`FJK3HSP_CP_R_QN_R, `FJK3HSP_CP_R_QN_F);
      if(IQ && CD && SD) (posedge CP => (QN +: K)) = (`FJK3HSP_CP_R_QN_R, `FJK3HSP_CP_R_QN_F);
      if(!SD) (posedge CD => (Q +: 1'b1)) = (`FJK3HSP_CD_R_Q_R,`FJK3HSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FJK3HSP_CD_R_Q_R,`FJK3HSP_CD_F_Q_F);
      if(CD) (negedge SD => (Q +: 1'b1)) = (`FJK3HSP_SD_F_Q_R,`FJK3HSP_SD_F_Q_R);
      if(!SD) (posedge CD => (QN +: 1'b0)) = (`FJK3HSP_CD_F_QN_R,`FJK3HSP_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`FJK3HSP_CD_F_QN_R,`FJK3HSP_CD_R_QN_F);
      if(CD) (negedge SD => (QN +: 1'b0)) = (`FJK3HSP_SD_F_QN_F,`FJK3HSP_SD_F_QN_F);

	$setuphold(posedge CP &&& AndCDSD_, posedge K, `FJK3HSP_K_CP_SETUP_posedge_posedge, `FJK3HSP_K_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSD_, negedge K, `FJK3HSP_K_CP_SETUP_negedge_posedge, `FJK3HSP_K_CP_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge CP &&& AndCDSD_, posedge J, `FJK3HSP_J_CP_SETUP_posedge_posedge, `FJK3HSP_J_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSD_, negedge J, `FJK3HSP_J_CP_SETUP_negedge_posedge, `FJK3HSP_J_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `FJK3HSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FJK3HSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FJK3HSP_SD_PWL, 0, Notifier);
      $width(negedge CD, `FJK3HSP_CD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& AndCDK, `FJK3HSP_SD_CP_REC_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge CP &&& AndSDJ, `FJK3HSP_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndCDK, posedge SD, `FJK3HSP_SD_CP_REM_posedge_posedge, Notifier);

	$hold(posedge CP &&& AndSDJ, posedge CD, `FJK3HSP_CD_CP_REM_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge SD, `FJK3HSP_CD_SD_REC_posedge_posedge, Notifier);

	$hold(posedge SD, posedge CD, `FJK3HSP_CD_SD_REM_posedge_posedge, Notifier);

`else

      (posedge CP => (Q +: Mux21JKXIQ_)) = (`FJK3HSP_CP_R_Q_R, `FJK3HSP_CP_R_Q_F);
      (posedge CP => (QN -: Mux21JKXIQ_)) = (`FJK3HSP_CP_R_QN_R, `FJK3HSP_CP_R_QN_F);
      (posedge CD => (Q +: 1'b1)) = (`FJK3HSP_CD_R_Q_R,`FJK3HSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`FJK3HSP_CD_R_Q_R,`FJK3HSP_CD_F_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`FJK3HSP_SD_F_Q_R,`FJK3HSP_SD_F_Q_R);
      (posedge CD => (QN +: 1'b0)) = (`FJK3HSP_CD_F_QN_R,`FJK3HSP_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`FJK3HSP_CD_F_QN_R,`FJK3HSP_CD_R_QN_F);
      (negedge SD => (QN +: 1'b0)) = (`FJK3HSP_SD_F_QN_F,`FJK3HSP_SD_F_QN_F);
 
        $setuphold(posedge CP &&& AndCDSD_, posedge K, `FJK3HSP_K_CP_SETUP_posedge_posedge, `FJK3HSP_K_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSD_, negedge K, `FJK3HSP_K_CP_SETUP_negedge_posedge, `FJK3HSP_K_CP_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge CP &&& AndCDSD_, posedge J, `FJK3HSP_J_CP_SETUP_posedge_posedge, `FJK3HSP_J_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSD_, negedge J, `FJK3HSP_J_CP_SETUP_negedge_posedge, `FJK3HSP_J_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `FJK3HSP_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `FJK3HSP_CP_PWH, 0, Notifier);
      $width(negedge SD, `FJK3HSP_SD_PWL, 0, Notifier);
      $width(negedge CD, `FJK3HSP_CD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& AndCDK, `FJK3HSP_SD_CP_REC_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge CP &&& AndSDJ, `FJK3HSP_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndCDK, posedge SD, `FJK3HSP_SD_CP_REM_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& AndSDJ, posedge CD, `FJK3HSP_CD_CP_REM_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge SD, `FJK3HSP_CD_SD_REC_posedge_posedge, Notifier);
 
        $hold(posedge SD, posedge CD, `FJK3HSP_CD_SD_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // FJK3HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:15 and Version :1.1 //
 
//  START 
// CELL HA01HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define HA01HS_B_F_CO_F 0.1
`define HA01HS_B_R_CO_R 0.1
`define HA01HS_A_F_CO_F 0.1
`define HA01HS_A_R_CO_R 0.1
`define HA01HS_B_F_S_R 0.1
`define HA01HS_B_R_S_F 0.1
`define HA01HS_B_F_S_F 0.1
`define HA01HS_B_R_S_R 0.1
`define HA01HS_A_F_S_R 0.1
`define HA01HS_A_R_S_F 0.1
`define HA01HS_A_F_S_F 0.1
`define HA01HS_A_R_S_R 0.1

module HA01HS (S, CO, A, B);

   output S;
   output CO;
   input A;
   input B;


   xor  u0 (S, A, B);
   and  u1 (CO, A, B);


`ifdef functional
`else
   specify

      (B +=> CO) = (`HA01HS_B_R_CO_R,`HA01HS_B_F_CO_F);
      (A +=> CO) = (`HA01HS_A_R_CO_R,`HA01HS_A_F_CO_F);
      if (A) (B -=> S) = (`HA01HS_B_F_S_R,`HA01HS_B_R_S_F);
      if (!A) (B +=> S) = (`HA01HS_B_R_S_R,`HA01HS_B_F_S_F);
      if (B) (A -=> S) = (`HA01HS_A_F_S_R,`HA01HS_A_R_S_F);
      if (!B) (A +=> S) = (`HA01HS_A_R_S_R,`HA01HS_A_F_S_F);

   endspecify
`endif


endmodule // HA01HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:26 and Version :1.1 //
 
// START
// CELL HA01HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define HA01HSP_B_F_CO_F 0.1
`define HA01HSP_B_R_CO_R 0.1
`define HA01HSP_A_F_CO_F 0.1
`define HA01HSP_A_R_CO_R 0.1
`define HA01HSP_B_F_S_R 0.1
`define HA01HSP_B_R_S_F 0.1
`define HA01HSP_B_F_S_F 0.1
`define HA01HSP_B_R_S_R 0.1
`define HA01HSP_A_F_S_R 0.1
`define HA01HSP_A_R_S_F 0.1
`define HA01HSP_A_F_S_F 0.1
`define HA01HSP_A_R_S_R 0.1

module HA01HSP (S, CO, A, B);

   output S;
   output CO;
   input A;
   input B;


   xor  u0 (S, A, B);
   and  u1 (CO, A, B);


`ifdef functional
`else
   specify

      (B +=> CO) = (`HA01HSP_B_R_CO_R,`HA01HSP_B_F_CO_F);
      (A +=> CO) = (`HA01HSP_A_R_CO_R,`HA01HSP_A_F_CO_F);
      if (A) (B -=> S) = (`HA01HSP_B_F_S_R,`HA01HSP_B_R_S_F);
      if (!A) (B +=> S) = (`HA01HSP_B_R_S_R,`HA01HSP_B_F_S_F);
      if (B) (A -=> S) = (`HA01HSP_A_F_S_R,`HA01HSP_A_R_S_F);
      if (!B) (A +=> S) = (`HA01HSP_A_R_S_R,`HA01HSP_A_F_S_F);

   endspecify
`endif


endmodule // HA01HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:26 and Version :1.1 //
 
// START
// CELL ITSHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ITSHS_E_F_Z_LZ 0.1
`define ITSHS_E_R_Z_ZL 0.1
`define ITSHS_E_F_Z_HZ 0.1
`define ITSHS_E_R_Z_ZH 0.1
`define ITSHS_A_F_Z_R 0.1
`define ITSHS_A_R_Z_F 0.1

module ITSHS (Z, A, E);

   output Z;
   input A;
   input E;


   notif1  u0 (Z, A, E);


`ifdef functional
`else
   specify

      (A -=> Z) = (`ITSHS_A_F_Z_R,`ITSHS_A_R_Z_F);
      (E => Z) = (`ITSHS_E_R_Z_ZH,`ITSHS_E_R_Z_ZL,`ITSHS_E_F_Z_LZ,`ITSHS_E_R_Z_ZH,`ITSHS_E_F_Z_HZ,`ITSHS_E_R_Z_ZL);

   endspecify
`endif


endmodule // ITSHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:29 and Version :1.1 //
 
//  START 
// CELL ITSHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ITSHSP_E_F_Z_LZ 0.1
`define ITSHSP_E_R_Z_ZL 0.1
`define ITSHSP_E_F_Z_HZ 0.1
`define ITSHSP_E_R_Z_ZH 0.1
`define ITSHSP_A_F_Z_R 0.1
`define ITSHSP_A_R_Z_F 0.1

module ITSHSP (Z, A, E);

   output Z;
   input A;
   input E;


   notif1  u0 (Z, A, E);


`ifdef functional
`else
   specify

      (A -=> Z) = (`ITSHSP_A_F_Z_R,`ITSHSP_A_R_Z_F);
      (E => Z) = (`ITSHSP_E_R_Z_ZH,`ITSHSP_E_R_Z_ZL,`ITSHSP_E_F_Z_LZ,`ITSHSP_E_R_Z_ZH,`ITSHSP_E_F_Z_HZ,`ITSHSP_E_R_Z_ZL);

   endspecify
`endif


endmodule // ITSHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:29 and Version :1.1 //
 
//  START 
// CELL ITSHSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ITSHSX3_E_F_Z_LZ 0.1
`define ITSHSX3_E_R_Z_ZL 0.1
`define ITSHSX3_E_F_Z_HZ 0.1
`define ITSHSX3_E_R_Z_ZH 0.1
`define ITSHSX3_A_F_Z_R 0.1
`define ITSHSX3_A_R_Z_F 0.1

module ITSHSX3 (Z, A, E);

   output Z;
   input A;
   input E;


   notif1  u0 (Z, A, E);


`ifdef functional
`else
   specify

      (A -=> Z) = (`ITSHSX3_A_F_Z_R,`ITSHSX3_A_R_Z_F);
      (E => Z) = (`ITSHSX3_E_R_Z_ZH,`ITSHSX3_E_R_Z_ZL,`ITSHSX3_E_F_Z_LZ,`ITSHSX3_E_R_Z_ZH,`ITSHSX3_E_F_Z_HZ,`ITSHSX3_E_R_Z_ZL);

   endspecify
`endif


endmodule // ITSHSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:29 and Version :1.1 //
 
//  START 
// CELL ITSHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ITSHSX4_E_F_Z_LZ 0.1
`define ITSHSX4_E_R_Z_ZL 0.1
`define ITSHSX4_E_F_Z_HZ 0.1
`define ITSHSX4_E_R_Z_ZH 0.1
`define ITSHSX4_A_F_Z_R 0.1
`define ITSHSX4_A_R_Z_F 0.1

module ITSHSX4 (Z, A, E);

   output Z;
   input A;
   input E;


   notif1  u0 (Z, A, E);


`ifdef functional
`else
   specify

      (A -=> Z) = (`ITSHSX4_A_F_Z_R,`ITSHSX4_A_R_Z_F);
      (E => Z) = (`ITSHSX4_E_R_Z_ZH,`ITSHSX4_E_R_Z_ZL,`ITSHSX4_E_F_Z_LZ,`ITSHSX4_E_R_Z_ZH,`ITSHSX4_E_F_Z_HZ,`ITSHSX4_E_R_Z_ZL);

   endspecify
`endif


endmodule // ITSHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:29 and Version :1.1 //
 
//  START 
// CELL ITSHSX5

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ITSHSX5_E_F_Z_LZ 0.1
`define ITSHSX5_E_R_Z_ZL 0.1
`define ITSHSX5_E_F_Z_HZ 0.1
`define ITSHSX5_E_R_Z_ZH 0.1
`define ITSHSX5_A_F_Z_R 0.1
`define ITSHSX5_A_R_Z_F 0.1

module ITSHSX5 (Z, A, E);

   output Z;
   input A;
   input E;


   notif1  u0 (Z, A, E);


`ifdef functional
`else
   specify

      (A -=> Z) = (`ITSHSX5_A_F_Z_R,`ITSHSX5_A_R_Z_F);
      (E => Z) = (`ITSHSX5_E_R_Z_ZH,`ITSHSX5_E_R_Z_ZL,`ITSHSX5_E_F_Z_LZ,`ITSHSX5_E_R_Z_ZH,`ITSHSX5_E_F_Z_HZ,`ITSHSX5_E_R_Z_ZL);

   endspecify
`endif


endmodule // ITSHSX5
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:29 and Version :1.1 //
 
//  START 
// CELL ITSHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ITSHSX8_E_F_Z_LZ 0.1
`define ITSHSX8_E_R_Z_ZL 0.1
`define ITSHSX8_E_F_Z_HZ 0.1
`define ITSHSX8_E_R_Z_ZH 0.1
`define ITSHSX8_A_F_Z_R 0.1
`define ITSHSX8_A_R_Z_F 0.1

module ITSHSX8 (Z, A, E);

   output Z;
   input A;
   input E;


   notif1  u0 (Z, A, E);


`ifdef functional
`else
   specify

      (A -=> Z) = (`ITSHSX8_A_F_Z_R,`ITSHSX8_A_R_Z_F);
      (E => Z) = (`ITSHSX8_E_R_Z_ZH,`ITSHSX8_E_R_Z_ZL,`ITSHSX8_E_F_Z_LZ,`ITSHSX8_E_R_Z_ZH,`ITSHSX8_E_F_Z_HZ,`ITSHSX8_E_R_Z_ZL);

   endspecify
`endif


endmodule // ITSHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:29 and Version :1.1 //
 
//  START 
// CELL ITSHSX16

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ITSHSX16_E_F_Z_LZ 0.1
`define ITSHSX16_E_R_Z_ZL 0.1
`define ITSHSX16_E_F_Z_HZ 0.1
`define ITSHSX16_E_R_Z_ZH 0.1
`define ITSHSX16_A_F_Z_R 0.1
`define ITSHSX16_A_R_Z_F 0.1

module ITSHSX16 (Z, A, E);

   output Z;
   input A;
   input E;


   notif1  u0 (Z, A, E);


`ifdef functional
`else
   specify

      (A -=> Z) = (`ITSHSX16_A_F_Z_R,`ITSHSX16_A_R_Z_F);
      (E => Z) = (`ITSHSX16_E_R_Z_ZH,`ITSHSX16_E_R_Z_ZL,`ITSHSX16_E_F_Z_LZ,`ITSHSX16_E_R_Z_ZH,`ITSHSX16_E_F_Z_HZ,`ITSHSX16_E_R_Z_ZL);

   endspecify
`endif


endmodule // ITSHSX16
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:29 and Version :1.1 //
 
//  START 
// CELL ITSHSX32

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ITSHSX32_E_F_Z_LZ 0.1
`define ITSHSX32_E_R_Z_ZL 0.1
`define ITSHSX32_E_F_Z_HZ 0.1
`define ITSHSX32_E_R_Z_ZH 0.1
`define ITSHSX32_A_F_Z_R 0.1
`define ITSHSX32_A_R_Z_F 0.1

module ITSHSX32 (Z, A, E);

   output Z;
   input A;
   input E;


   notif1  u0 (Z, A, E);


`ifdef functional
`else
   specify

      (A -=> Z) = (`ITSHSX32_A_F_Z_R,`ITSHSX32_A_R_Z_F);
      (E => Z) = (`ITSHSX32_E_R_Z_ZH,`ITSHSX32_E_R_Z_ZL,`ITSHSX32_E_F_Z_LZ,`ITSHSX32_E_R_Z_ZH,`ITSHSX32_E_F_Z_HZ,`ITSHSX32_E_R_Z_ZL);

   endspecify
`endif


endmodule // ITSHSX32
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:29 and Version :1.1 //
 
//  START 
// CELL ITSENHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ITSENHS_EN_F_Z_ZL 0.1
`define ITSENHS_EN_R_Z_LZ 0.1
`define ITSENHS_EN_F_Z_ZH 0.1
`define ITSENHS_EN_R_Z_HZ 0.1
`define ITSENHS_A_F_Z_R 0.1
`define ITSENHS_A_R_Z_F 0.1

module ITSENHS (Z, A, EN);

   output Z;
   input A;
   input EN;


   notif0  u0 (Z, A, EN);


`ifdef functional
`else
   specify

      (A -=> Z) = (`ITSENHS_A_F_Z_R,`ITSENHS_A_R_Z_F);
      (EN => Z) = (`ITSENHS_EN_F_Z_ZH,`ITSENHS_EN_F_Z_ZL,`ITSENHS_EN_R_Z_LZ,`ITSENHS_EN_F_Z_ZH,`ITSENHS_EN_R_Z_HZ,`ITSENHS_EN_F_Z_ZL);

   endspecify
`endif


endmodule // ITSENHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:29 and Version :1.1 //
 
//  START 
// CELL ITSENHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ITSENHSP_EN_F_Z_ZL 0.1
`define ITSENHSP_EN_R_Z_LZ 0.1
`define ITSENHSP_EN_F_Z_ZH 0.1
`define ITSENHSP_EN_R_Z_HZ 0.1
`define ITSENHSP_A_F_Z_R 0.1
`define ITSENHSP_A_R_Z_F 0.1

module ITSENHSP (Z, A, EN);

   output Z;
   input A;
   input EN;


   notif0  u0 (Z, A, EN);


`ifdef functional
`else
   specify

      (A -=> Z) = (`ITSENHSP_A_F_Z_R,`ITSENHSP_A_R_Z_F);
      (EN => Z) = (`ITSENHSP_EN_F_Z_ZH,`ITSENHSP_EN_F_Z_ZL,`ITSENHSP_EN_R_Z_LZ,`ITSENHSP_EN_F_Z_ZH,`ITSENHSP_EN_R_Z_HZ,`ITSENHSP_EN_F_Z_ZL);

   endspecify
`endif


endmodule // ITSENHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:29 and Version :1.1 //
 
//  START 
// CELL ITSENHSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ITSENHSX3_EN_F_Z_ZL 0.1
`define ITSENHSX3_EN_R_Z_LZ 0.1
`define ITSENHSX3_EN_F_Z_ZH 0.1
`define ITSENHSX3_EN_R_Z_HZ 0.1
`define ITSENHSX3_A_F_Z_R 0.1
`define ITSENHSX3_A_R_Z_F 0.1

module ITSENHSX3 (Z, A, EN);

   output Z;
   input A;
   input EN;


   notif0  u0 (Z, A, EN);


`ifdef functional
`else
   specify

      (A -=> Z) = (`ITSENHSX3_A_F_Z_R,`ITSENHSX3_A_R_Z_F);
      (EN => Z) = (`ITSENHSX3_EN_F_Z_ZH,`ITSENHSX3_EN_F_Z_ZL,`ITSENHSX3_EN_R_Z_LZ,`ITSENHSX3_EN_F_Z_ZH,`ITSENHSX3_EN_R_Z_HZ,`ITSENHSX3_EN_F_Z_ZL);

   endspecify
`endif


endmodule // ITSENHSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:29 and Version :1.1 //
 
//  START 
// CELL ITSENHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ITSENHSX4_EN_F_Z_ZL 0.1
`define ITSENHSX4_EN_R_Z_LZ 0.1
`define ITSENHSX4_EN_F_Z_ZH 0.1
`define ITSENHSX4_EN_R_Z_HZ 0.1
`define ITSENHSX4_A_F_Z_R 0.1
`define ITSENHSX4_A_R_Z_F 0.1

module ITSENHSX4 (Z, A, EN);

   output Z;
   input A;
   input EN;


   notif0  u0 (Z, A, EN);


`ifdef functional
`else
   specify

      (A -=> Z) = (`ITSENHSX4_A_F_Z_R,`ITSENHSX4_A_R_Z_F);
      (EN => Z) = (`ITSENHSX4_EN_F_Z_ZH,`ITSENHSX4_EN_F_Z_ZL,`ITSENHSX4_EN_R_Z_LZ,`ITSENHSX4_EN_F_Z_ZH,`ITSENHSX4_EN_R_Z_HZ,`ITSENHSX4_EN_F_Z_ZL);

   endspecify
`endif


endmodule // ITSENHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:29 and Version :1.1 //
 
//  START 
// CELL ITSENHSX5

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ITSENHSX5_EN_F_Z_ZL 0.1
`define ITSENHSX5_EN_R_Z_LZ 0.1
`define ITSENHSX5_EN_F_Z_ZH 0.1
`define ITSENHSX5_EN_R_Z_HZ 0.1
`define ITSENHSX5_A_F_Z_R 0.1
`define ITSENHSX5_A_R_Z_F 0.1

module ITSENHSX5 (Z, A, EN);

   output Z;
   input A;
   input EN;


   notif0  u0 (Z, A, EN);


`ifdef functional
`else
   specify

      (A -=> Z) = (`ITSENHSX5_A_F_Z_R,`ITSENHSX5_A_R_Z_F);
      (EN => Z) = (`ITSENHSX5_EN_F_Z_ZH,`ITSENHSX5_EN_F_Z_ZL,`ITSENHSX5_EN_R_Z_LZ,`ITSENHSX5_EN_F_Z_ZH,`ITSENHSX5_EN_R_Z_HZ,`ITSENHSX5_EN_F_Z_ZL);

   endspecify
`endif


endmodule // ITSENHSX5
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:29 and Version :1.1 //
 
//  START 
// CELL ITSENHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ITSENHSX8_EN_F_Z_ZL 0.1
`define ITSENHSX8_EN_R_Z_LZ 0.1
`define ITSENHSX8_EN_F_Z_ZH 0.1
`define ITSENHSX8_EN_R_Z_HZ 0.1
`define ITSENHSX8_A_F_Z_R 0.1
`define ITSENHSX8_A_R_Z_F 0.1

module ITSENHSX8 (Z, A, EN);

   output Z;
   input A;
   input EN;


   notif0  u0 (Z, A, EN);


`ifdef functional
`else
   specify

      (A -=> Z) = (`ITSENHSX8_A_F_Z_R,`ITSENHSX8_A_R_Z_F);
      (EN => Z) = (`ITSENHSX8_EN_F_Z_ZH,`ITSENHSX8_EN_F_Z_ZL,`ITSENHSX8_EN_R_Z_LZ,`ITSENHSX8_EN_F_Z_ZH,`ITSENHSX8_EN_R_Z_HZ,`ITSENHSX8_EN_F_Z_ZL);

   endspecify
`endif


endmodule // ITSENHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:29 and Version :1.1 //
 
//  START 
// CELL ITSENHSX16

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ITSENHSX16_EN_F_Z_ZL 0.1
`define ITSENHSX16_EN_R_Z_LZ 0.1
`define ITSENHSX16_EN_F_Z_ZH 0.1
`define ITSENHSX16_EN_R_Z_HZ 0.1
`define ITSENHSX16_A_F_Z_R 0.1
`define ITSENHSX16_A_R_Z_F 0.1

module ITSENHSX16 (Z, A, EN);

   output Z;
   input A;
   input EN;


   notif0  u0 (Z, A, EN);


`ifdef functional
`else
   specify

      (A -=> Z) = (`ITSENHSX16_A_F_Z_R,`ITSENHSX16_A_R_Z_F);
      (EN => Z) = (`ITSENHSX16_EN_F_Z_ZH,`ITSENHSX16_EN_F_Z_ZL,`ITSENHSX16_EN_R_Z_LZ,`ITSENHSX16_EN_F_Z_ZH,`ITSENHSX16_EN_R_Z_HZ,`ITSENHSX16_EN_F_Z_ZL);

   endspecify
`endif


endmodule // ITSENHSX16
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:29 and Version :1.1 //
 
//  START 
// CELL ITSENHSX32

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ITSENHSX32_EN_F_Z_ZL 0.1
`define ITSENHSX32_EN_R_Z_LZ 0.1
`define ITSENHSX32_EN_F_Z_ZH 0.1
`define ITSENHSX32_EN_R_Z_HZ 0.1
`define ITSENHSX32_A_F_Z_R 0.1
`define ITSENHSX32_A_R_Z_F 0.1

module ITSENHSX32 (Z, A, EN);

   output Z;
   input A;
   input EN;


   notif0  u0 (Z, A, EN);


`ifdef functional
`else
   specify

      (A -=> Z) = (`ITSENHSX32_A_F_Z_R,`ITSENHSX32_A_R_Z_F);
      (EN => Z) = (`ITSENHSX32_EN_F_Z_ZH,`ITSENHSX32_EN_F_Z_ZL,`ITSENHSX32_EN_R_Z_LZ,`ITSENHSX32_EN_F_Z_ZH,`ITSENHSX32_EN_R_Z_HZ,`ITSENHSX32_EN_F_Z_ZL);

   endspecify
`endif


endmodule // ITSENHSX32
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:29 and Version :1.1 //
 
//  START 
// CELL IVHSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define IVHSX05_A_F_Z_R 0.1
`define IVHSX05_A_R_Z_F 0.1

module IVHSX05 (Z, A);

   output Z;
   input A;


   not  u0 (Z, A);


`ifdef functional
`else
   specify

      (A -=> Z) = (`IVHSX05_A_F_Z_R,`IVHSX05_A_R_Z_F);

   endspecify
`endif


endmodule // IVHSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:33 and Version :1.1 //
 
//  START
// CELL IVHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define IVHS_A_F_Z_R 0.1
`define IVHS_A_R_Z_F 0.1

module IVHS (Z, A);

   output Z;
   input A;


   not  u0 (Z, A);


`ifdef functional
`else
   specify

      (A -=> Z) = (`IVHS_A_F_Z_R,`IVHS_A_R_Z_F);

   endspecify
`endif


endmodule // IVHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:33 and Version :1.1 //
 
//  START
// CELL IVHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define IVHSP_A_F_Z_R 0.1
`define IVHSP_A_R_Z_F 0.1

module IVHSP (Z, A);

   output Z;
   input A;


   not  u0 (Z, A);


`ifdef functional
`else
   specify

      (A -=> Z) = (`IVHSP_A_F_Z_R,`IVHSP_A_R_Z_F);

   endspecify
`endif


endmodule // IVHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:33 and Version :1.1 //
 
//  START
// CELL IVHSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define IVHSX3_A_F_Z_R 0.1
`define IVHSX3_A_R_Z_F 0.1

module IVHSX3 (Z, A);

   output Z;
   input A;


   not  u0 (Z, A);


`ifdef functional
`else
   specify

      (A -=> Z) = (`IVHSX3_A_F_Z_R,`IVHSX3_A_R_Z_F);

   endspecify
`endif


endmodule // IVHSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:33 and Version :1.1 //
 
//  START
// CELL IVHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define IVHSX4_A_F_Z_R 0.1
`define IVHSX4_A_R_Z_F 0.1

module IVHSX4 (Z, A);

   output Z;
   input A;


   not  u0 (Z, A);


`ifdef functional
`else
   specify

      (A -=> Z) = (`IVHSX4_A_F_Z_R,`IVHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // IVHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:33 and Version :1.1 //
 
//  START
// CELL IVHSX5

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define IVHSX5_A_F_Z_R 0.1
`define IVHSX5_A_R_Z_F 0.1

module IVHSX5 (Z, A);

   output Z;
   input A;


   not  u0 (Z, A);


`ifdef functional
`else
   specify

      (A -=> Z) = (`IVHSX5_A_F_Z_R,`IVHSX5_A_R_Z_F);

   endspecify
`endif


endmodule // IVHSX5
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:33 and Version :1.1 //
 
//  START
// CELL IVHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define IVHSX8_A_F_Z_R 0.1
`define IVHSX8_A_R_Z_F 0.1

module IVHSX8 (Z, A);

   output Z;
   input A;


   not  u0 (Z, A);


`ifdef functional
`else
   specify

      (A -=> Z) = (`IVHSX8_A_F_Z_R,`IVHSX8_A_R_Z_F);

   endspecify
`endif


endmodule // IVHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:33 and Version :1.1 //
 
//  START
// CELL IVHSX16

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define IVHSX16_A_F_Z_R 0.1
`define IVHSX16_A_R_Z_F 0.1

module IVHSX16 (Z, A);

   output Z;
   input A;


   not  u0 (Z, A);


`ifdef functional
`else
   specify

      (A -=> Z) = (`IVHSX16_A_F_Z_R,`IVHSX16_A_R_Z_F);

   endspecify
`endif


endmodule // IVHSX16
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:33 and Version :1.1 //
 
//  START
// CELL IVHSX32

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define IVHSX32_A_F_Z_R 0.1
`define IVHSX32_A_R_Z_F 0.1

module IVHSX32 (Z, A);

   output Z;
   input A;


   not  u0 (Z, A);


`ifdef functional
`else
   specify

      (A -=> Z) = (`IVHSX32_A_F_Z_R,`IVHSX32_A_R_Z_F);

   endspecify
`endif


endmodule // IVHSX32
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:33 and Version :1.1 //
 
//  START
// CELL F_IVHSX16

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_IVHSX16_A_F_Z_R 0.1
`define F_IVHSX16_A_R_Z_F 0.1

module F_IVHSX16 (Z, A);

   output Z;
   input A;


   not  u0 (Z, A);


`ifdef functional
`else
   specify

      (A -=> Z) = (`F_IVHSX16_A_F_Z_R,`F_IVHSX16_A_R_Z_F);

   endspecify
`endif


endmodule // F_IVHSX16
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:33 and Version :1.1 //
 
//  START
// CELL F_IVHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_IVHSX8_A_F_Z_R 0.1
`define F_IVHSX8_A_R_Z_F 0.1

module F_IVHSX8 (Z, A);

   output Z;
   input A;


   not  u0 (Z, A);


`ifdef functional
`else
   specify

      (A -=> Z) = (`F_IVHSX8_A_F_Z_R,`F_IVHSX8_A_R_Z_F);

   endspecify
`endif


endmodule // F_IVHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:33 and Version :1.1 //
 
//  START
// CELL M_IVHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define M_IVHSP_A_F_Z_R 0.1
`define M_IVHSP_A_R_Z_F 0.1

module M_IVHSP (Z, A);

   output Z;
   input A;


   not  u0 (Z, A);


`ifdef functional
`else
   specify

      (A -=> Z) = (`M_IVHSP_A_F_Z_R,`M_IVHSP_A_R_Z_F);

   endspecify
`endif


endmodule // M_IVHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:33 and Version :1.1 //
 
//  START
// CELL M_IVHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define M_IVHSX4_A_F_Z_R 0.1
`define M_IVHSX4_A_R_Z_F 0.1

module M_IVHSX4 (Z, A);

   output Z;
   input A;


   not  u0 (Z, A);


`ifdef functional
`else
   specify

      (A -=> Z) = (`M_IVHSX4_A_F_Z_R,`M_IVHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // M_IVHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:33 and Version :1.1 //
 
//  START
// CELL LD1HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD1HS_G_R_QN_F 0.1
`define LD1HS_G_R_QN_R 0.1
`define LD1HS_D_F_QN_R 0.1
`define LD1HS_D_R_QN_F 0.1
`define LD1HS_G_R_Q_R 0.1
`define LD1HS_G_R_Q_F 0.1
`define LD1HS_D_F_Q_F 0.1
`define LD1HS_D_R_Q_R 0.1
`define LD1HS_G_PWH 0.1
`define LD1HS_D_G_SETUP_posedge_negedge 0.1
`define LD1HS_D_G_SETUP_negedge_negedge 0.1
`define LD1HS_D_G_HOLD_posedge_negedge 0.1
`define LD1HS_D_G_HOLD_negedge_negedge 0.1

module LD1HS (Q, QN, D, G);

   output Q;
   output QN;
   input D;
   input G;


   reg Notifier;


   U_LD_P_NOTI u0 (   // Verilog Seq UDP
      IQ, D, G, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   specify

      if (G) (D -=> QN) = (`LD1HS_D_F_QN_R,`LD1HS_D_R_QN_F);
      if (G) (D +=> Q) = (`LD1HS_D_R_Q_R,`LD1HS_D_F_Q_F);
      (posedge G => (Q +: D)) = (`LD1HS_G_R_Q_R, `LD1HS_G_R_Q_F);
      (posedge G => (QN -: D)) = (`LD1HS_G_R_QN_R, `LD1HS_G_R_QN_F);

	$setuphold(negedge G, posedge D, `LD1HS_D_G_SETUP_posedge_negedge, `LD1HS_D_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G, negedge D, `LD1HS_D_G_SETUP_negedge_negedge, `LD1HS_D_G_HOLD_negedge_negedge, Notifier);

      $width(posedge G, `LD1HS_G_PWH, 0, Notifier);

   endspecify
`endif


endmodule // LD1HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:35 and Version :1.1 //
 
//  START 
// CELL LD1HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD1HSP_G_R_QN_F 0.1
`define LD1HSP_G_R_QN_R 0.1
`define LD1HSP_D_F_QN_R 0.1
`define LD1HSP_D_R_QN_F 0.1
`define LD1HSP_G_R_Q_R 0.1
`define LD1HSP_G_R_Q_F 0.1
`define LD1HSP_D_F_Q_F 0.1
`define LD1HSP_D_R_Q_R 0.1
`define LD1HSP_G_PWH 0.1
`define LD1HSP_D_G_SETUP_posedge_negedge 0.1
`define LD1HSP_D_G_SETUP_negedge_negedge 0.1
`define LD1HSP_D_G_HOLD_posedge_negedge 0.1
`define LD1HSP_D_G_HOLD_negedge_negedge 0.1

module LD1HSP (Q, QN, D, G);

   output Q;
   output QN;
   input D;
   input G;


   reg Notifier;


   U_LD_P_NOTI u0 (   // Verilog Seq UDP
      IQ, D, G, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   specify

      if (G) (D -=> QN) = (`LD1HSP_D_F_QN_R,`LD1HSP_D_R_QN_F);
      if (G) (D +=> Q) = (`LD1HSP_D_R_Q_R,`LD1HSP_D_F_Q_F);
      (posedge G => (Q +: D)) = (`LD1HSP_G_R_Q_R, `LD1HSP_G_R_Q_F);
      (posedge G => (QN -: D)) = (`LD1HSP_G_R_QN_R, `LD1HSP_G_R_QN_F);

	$setuphold(negedge G, posedge D, `LD1HSP_D_G_SETUP_posedge_negedge, `LD1HSP_D_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G, negedge D, `LD1HSP_D_G_SETUP_negedge_negedge, `LD1HSP_D_G_HOLD_negedge_negedge, Notifier);

      $width(posedge G, `LD1HSP_G_PWH, 0, Notifier);

   endspecify
`endif


endmodule // LD1HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:35 and Version :1.1 //
 
//  START 
// CELL LD1QHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD1QHS_G_R_Q_R 0.1
`define LD1QHS_G_R_Q_F 0.1
`define LD1QHS_D_F_Q_F 0.1
`define LD1QHS_D_R_Q_R 0.1
`define LD1QHS_D_G_HOLD_posedge_negedge 0.1
`define LD1QHS_D_G_HOLD_negedge_negedge 0.1
`define LD1QHS_D_G_SETUP_posedge_negedge 0.1
`define LD1QHS_D_G_SETUP_negedge_negedge 0.1
`define LD1QHS_G_PWH 0.1

module LD1QHS (Q, D, G);

   output Q;
   input D;
   input G;


   reg Notifier;


   U_LD_P_NOTI u0 (IQ, D, G, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify

      if (G) (D +=> Q) = (`LD1QHS_D_R_Q_R,`LD1QHS_D_F_Q_F);
      (posedge G => (Q +: D)) = (`LD1QHS_G_R_Q_R, `LD1QHS_G_R_Q_F);

	$setuphold(negedge G, posedge D, `LD1QHS_D_G_SETUP_posedge_negedge, `LD1QHS_D_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G, negedge D, `LD1QHS_D_G_SETUP_negedge_negedge, `LD1QHS_D_G_HOLD_negedge_negedge, Notifier);

      $width(posedge G, `LD1QHS_G_PWH, 0, Notifier);

   endspecify
`endif


endmodule // LD1QHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:39 and Version :1.1 //
 
//  START 
// CELL LD1QHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD1QHSP_G_R_Q_R 0.1
`define LD1QHSP_G_R_Q_F 0.1
`define LD1QHSP_D_F_Q_F 0.1
`define LD1QHSP_D_R_Q_R 0.1
`define LD1QHSP_D_G_HOLD_posedge_negedge 0.1
`define LD1QHSP_D_G_HOLD_negedge_negedge 0.1
`define LD1QHSP_D_G_SETUP_posedge_negedge 0.1
`define LD1QHSP_D_G_SETUP_negedge_negedge 0.1
`define LD1QHSP_G_PWH 0.1

module LD1QHSP (Q, D, G);

   output Q;
   input D;
   input G;


   reg Notifier;


   U_LD_P_NOTI u0 (IQ, D, G, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify

      if (G) (D +=> Q) = (`LD1QHSP_D_R_Q_R,`LD1QHSP_D_F_Q_F);
      (posedge G => (Q +: D)) = (`LD1QHSP_G_R_Q_R, `LD1QHSP_G_R_Q_F);

	$setuphold(negedge G, posedge D, `LD1QHSP_D_G_SETUP_posedge_negedge, `LD1QHSP_D_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G, negedge D, `LD1QHSP_D_G_SETUP_negedge_negedge, `LD1QHSP_D_G_HOLD_negedge_negedge, Notifier);

      $width(posedge G, `LD1QHSP_G_PWH, 0, Notifier);

   endspecify
`endif


endmodule // LD1QHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:39 and Version :1.1 //
 
//  START 
// CELL LD1QHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD1QHSX4_G_R_Q_R 0.1
`define LD1QHSX4_G_R_Q_F 0.1
`define LD1QHSX4_D_F_Q_F 0.1
`define LD1QHSX4_D_R_Q_R 0.1
`define LD1QHSX4_D_G_HOLD_posedge_negedge 0.1
`define LD1QHSX4_D_G_HOLD_negedge_negedge 0.1
`define LD1QHSX4_D_G_SETUP_posedge_negedge 0.1
`define LD1QHSX4_D_G_SETUP_negedge_negedge 0.1
`define LD1QHSX4_G_PWH 0.1

module LD1QHSX4 (Q, D, G);

   output Q;
   input D;
   input G;


   reg Notifier;


   U_LD_P_NOTI u0 (IQ, D, G, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify

      if (G) (D +=> Q) = (`LD1QHSX4_D_R_Q_R,`LD1QHSX4_D_F_Q_F);
      (posedge G => (Q +: D)) = (`LD1QHSX4_G_R_Q_R, `LD1QHSX4_G_R_Q_F);

	$setuphold(negedge G, posedge D, `LD1QHSX4_D_G_SETUP_posedge_negedge, `LD1QHSX4_D_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G, negedge D, `LD1QHSX4_D_G_SETUP_negedge_negedge, `LD1QHSX4_D_G_HOLD_negedge_negedge, Notifier);

      $width(posedge G, `LD1QHSX4_G_PWH, 0, Notifier);

   endspecify
`endif


endmodule // LD1QHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:39 and Version :1.1 //
 
//  START 
// CELL LD1SHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD1SHS_TE_F_QN_R 0.1
`define LD1SHS_TE_R_QN_F 0.1
`define LD1SHS_TE_F_QN_F 0.1
`define LD1SHS_TE_R_QN_R 0.1
`define LD1SHS_TI_F_QN_R 0.1
`define LD1SHS_TI_R_QN_F 0.1
`define LD1SHS_G_R_QN_F 0.1
`define LD1SHS_G_R_QN_R 0.1
`define LD1SHS_D_F_QN_R 0.1
`define LD1SHS_D_R_QN_F 0.1
`define LD1SHS_TE_F_Q_F 0.1
`define LD1SHS_TE_R_Q_R 0.1
`define LD1SHS_TE_F_Q_R 0.1
`define LD1SHS_TE_R_Q_F 0.1
`define LD1SHS_TI_F_Q_F 0.1
`define LD1SHS_TI_R_Q_R 0.1
`define LD1SHS_G_R_Q_R 0.1
`define LD1SHS_G_R_Q_F 0.1
`define LD1SHS_D_F_Q_F 0.1
`define LD1SHS_D_R_Q_R 0.1
`define LD1SHS_G_PWH 0.1
`define LD1SHS_D_G_SETUP_posedge_negedge 0.1
`define LD1SHS_D_G_SETUP_negedge_negedge 0.1
`define LD1SHS_D_G_HOLD_posedge_negedge 0.1
`define LD1SHS_D_G_HOLD_negedge_negedge 0.1
`define LD1SHS_TI_G_SETUP_posedge_negedge 0.1
`define LD1SHS_TI_G_SETUP_negedge_negedge 0.1
`define LD1SHS_TI_G_HOLD_posedge_negedge 0.1
`define LD1SHS_TI_G_HOLD_negedge_negedge 0.1
`define LD1SHS_TE_G_SETUP_posedge_negedge 0.1
`define LD1SHS_TE_G_SETUP_negedge_negedge 0.1
`define LD1SHS_TE_G_HOLD_posedge_negedge 0.1
`define LD1SHS_TE_G_HOLD_negedge_negedge 0.1

module LD1SHS (Q, QN, D, G, TI, TE);

   output Q;
   output QN;
   input D;
   input G;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_LD_P_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, G, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault
 
      if (!D && G && TI) (TE -=> QN) = (`LD1SHS_TE_F_QN_R,`LD1SHS_TE_R_QN_F);
      if (D && G && !TI) (TE +=> QN) = (`LD1SHS_TE_R_QN_R,`LD1SHS_TE_F_QN_F);
      if (G && TE) (TI -=> QN) = (`LD1SHS_TI_F_QN_R,`LD1SHS_TI_R_QN_F);
      if (G && !TE) (D -=> QN) = (`LD1SHS_D_F_QN_R,`LD1SHS_D_R_QN_F);
      if (!D && G && TI) (TE +=> Q) = (`LD1SHS_TE_R_Q_R,`LD1SHS_TE_F_Q_F);
      if (D && G && !TI) (TE -=> Q) = (`LD1SHS_TE_F_Q_R,`LD1SHS_TE_R_Q_F);
      if (G && TE) (TI +=> Q) = (`LD1SHS_TI_R_Q_R,`LD1SHS_TI_F_Q_F);
      if (G && !TE) (D +=> Q) = (`LD1SHS_D_R_Q_R,`LD1SHS_D_F_Q_F);
      if(!TE) (posedge G => (Q +: D)) = (`LD1SHS_G_R_Q_R, `LD1SHS_G_R_Q_F);
      if(TE) (posedge G => (Q +: TI)) = (`LD1SHS_G_R_Q_R, `LD1SHS_G_R_Q_F);
      if(!D && TI) (posedge G => (Q +: TE)) = (`LD1SHS_G_R_Q_R, `LD1SHS_G_R_Q_F);
      if(!TI && D) (posedge G => (Q -: TE)) = (`LD1SHS_G_R_Q_R, `LD1SHS_G_R_Q_F);
      if(!TE) (posedge G => (QN -: D)) = (`LD1SHS_G_R_QN_R, `LD1SHS_G_R_QN_F);
      if(TE) (posedge G => (QN -: TI)) = (`LD1SHS_G_R_QN_R, `LD1SHS_G_R_QN_F);
      if(!D && TI) (posedge G => (QN -: TE)) = (`LD1SHS_G_R_QN_R, `LD1SHS_G_R_QN_F);
      if(!TI && D) (posedge G => (QN +: TE)) = (`LD1SHS_G_R_QN_R, `LD1SHS_G_R_QN_F);

	$setuphold(negedge G &&& XorDTI_, posedge TE, `LD1SHS_TE_G_SETUP_posedge_negedge, `LD1SHS_TE_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& XorDTI_, negedge TE, `LD1SHS_TE_G_SETUP_negedge_negedge, `LD1SHS_TE_G_HOLD_negedge_negedge, Notifier);

	$setuphold(negedge G &&& TE, posedge TI, `LD1SHS_TI_G_SETUP_posedge_negedge, `LD1SHS_TI_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& TE, negedge TI, `LD1SHS_TI_G_SETUP_negedge_negedge, `LD1SHS_TI_G_HOLD_negedge_negedge, Notifier);

	$setuphold(negedge G &&& TEX, posedge D, `LD1SHS_D_G_SETUP_posedge_negedge, `LD1SHS_D_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& TEX, negedge D, `LD1SHS_D_G_SETUP_negedge_negedge, `LD1SHS_D_G_HOLD_negedge_negedge, Notifier);

      $width(posedge G, `LD1SHS_G_PWH, 0, Notifier);
`else

     if (!D && G && TI) (TE -=> QN) = (`LD1SHS_TE_F_QN_R,`LD1SHS_TE_R_QN_F);
     if (D && G && !TI) (TE +=> QN) = (`LD1SHS_TE_R_QN_R,`LD1SHS_TE_F_QN_F);
      (TI -=> QN) = (`LD1SHS_TI_F_QN_R,`LD1SHS_TI_R_QN_F);
      (D -=> QN) = (`LD1SHS_D_F_QN_R,`LD1SHS_D_R_QN_F);
     if (!D && G && TI) (TE +=> Q) = (`LD1SHS_TE_R_Q_R,`LD1SHS_TE_F_Q_F);
      if (D && G && !TI) (TE -=> Q) = (`LD1SHS_TE_F_Q_R,`LD1SHS_TE_R_Q_F);
      (TI +=> Q) = (`LD1SHS_TI_R_Q_R,`LD1SHS_TI_F_Q_F);
      (D +=> Q) = (`LD1SHS_D_R_Q_R,`LD1SHS_D_F_Q_F);
      (posedge G => (Q +: Mux21DTITE_)) = (`LD1SHS_G_R_Q_R, `LD1SHS_G_R_Q_F);
      (posedge G => (QN -: Mux21DTITE_)) = (`LD1SHS_G_R_QN_R, `LD1SHS_G_R_QN_F);
 
        $setuphold(negedge G &&& XorDTI_, posedge TE, `LD1SHS_TE_G_SETUP_posedge_negedge, `LD1SHS_TE_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& XorDTI_, negedge TE, `LD1SHS_TE_G_SETUP_negedge_negedge, `LD1SHS_TE_G_HOLD_negedge_negedge, Notifier);
 
        $setuphold(negedge G &&& TE, posedge TI, `LD1SHS_TI_G_SETUP_posedge_negedge, `LD1SHS_TI_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& TE, negedge TI, `LD1SHS_TI_G_SETUP_negedge_negedge, `LD1SHS_TI_G_HOLD_negedge_negedge, Notifier);
 
        $setuphold(negedge G &&& TEX, posedge D, `LD1SHS_D_G_SETUP_posedge_negedge, `LD1SHS_D_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& TEX, negedge D, `LD1SHS_D_G_SETUP_negedge_negedge, `LD1SHS_D_G_HOLD_negedge_negedge, Notifier);
 
      $width(posedge G, `LD1SHS_G_PWH, 0, Notifier);
`endif
   endspecify
`endif


endmodule // LD1SHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:45 and Version :1.1 //
 
//  START 
// CELL LD1SHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD1SHSP_TE_F_QN_R 0.1
`define LD1SHSP_TE_R_QN_F 0.1
`define LD1SHSP_TE_F_QN_F 0.1
`define LD1SHSP_TE_R_QN_R 0.1
`define LD1SHSP_TI_F_QN_R 0.1
`define LD1SHSP_TI_R_QN_F 0.1
`define LD1SHSP_G_R_QN_F 0.1
`define LD1SHSP_G_R_QN_R 0.1
`define LD1SHSP_D_F_QN_R 0.1
`define LD1SHSP_D_R_QN_F 0.1
`define LD1SHSP_TE_F_Q_F 0.1
`define LD1SHSP_TE_R_Q_R 0.1
`define LD1SHSP_TE_F_Q_R 0.1
`define LD1SHSP_TE_R_Q_F 0.1
`define LD1SHSP_TI_F_Q_F 0.1
`define LD1SHSP_TI_R_Q_R 0.1
`define LD1SHSP_G_R_Q_R 0.1
`define LD1SHSP_G_R_Q_F 0.1
`define LD1SHSP_D_F_Q_F 0.1
`define LD1SHSP_D_R_Q_R 0.1
`define LD1SHSP_G_PWH 0.1
`define LD1SHSP_D_G_SETUP_posedge_negedge 0.1
`define LD1SHSP_D_G_SETUP_negedge_negedge 0.1
`define LD1SHSP_D_G_HOLD_posedge_negedge 0.1
`define LD1SHSP_D_G_HOLD_negedge_negedge 0.1
`define LD1SHSP_TI_G_SETUP_posedge_negedge 0.1
`define LD1SHSP_TI_G_SETUP_negedge_negedge 0.1
`define LD1SHSP_TI_G_HOLD_posedge_negedge 0.1
`define LD1SHSP_TI_G_HOLD_negedge_negedge 0.1
`define LD1SHSP_TE_G_SETUP_posedge_negedge 0.1
`define LD1SHSP_TE_G_SETUP_negedge_negedge 0.1
`define LD1SHSP_TE_G_HOLD_posedge_negedge 0.1
`define LD1SHSP_TE_G_HOLD_negedge_negedge 0.1

module LD1SHSP (Q, QN, D, G, TI, TE);

   output Q;
   output QN;
   input D;
   input G;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_LD_P_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, G, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault
 
      if (!D && G && TI) (TE -=> QN) = (`LD1SHSP_TE_F_QN_R,`LD1SHSP_TE_R_QN_F);
      if (D && G && !TI) (TE +=> QN) = (`LD1SHSP_TE_R_QN_R,`LD1SHSP_TE_F_QN_F);
      if (G && TE) (TI -=> QN) = (`LD1SHSP_TI_F_QN_R,`LD1SHSP_TI_R_QN_F);
      if (G && !TE) (D -=> QN) = (`LD1SHSP_D_F_QN_R,`LD1SHSP_D_R_QN_F);
      if (!D && G && TI) (TE +=> Q) = (`LD1SHSP_TE_R_Q_R,`LD1SHSP_TE_F_Q_F);
      if (D && G && !TI) (TE -=> Q) = (`LD1SHSP_TE_F_Q_R,`LD1SHSP_TE_R_Q_F);
      if (G && TE) (TI +=> Q) = (`LD1SHSP_TI_R_Q_R,`LD1SHSP_TI_F_Q_F);
      if (G && !TE) (D +=> Q) = (`LD1SHSP_D_R_Q_R,`LD1SHSP_D_F_Q_F);
      if(!TE) (posedge G => (Q +: D)) = (`LD1SHSP_G_R_Q_R, `LD1SHSP_G_R_Q_F);
      if(TE) (posedge G => (Q +: TI)) = (`LD1SHSP_G_R_Q_R, `LD1SHSP_G_R_Q_F);
      if(!D && TI) (posedge G => (Q +: TE)) = (`LD1SHSP_G_R_Q_R, `LD1SHSP_G_R_Q_F);
      if(!TI && D) (posedge G => (Q -: TE)) = (`LD1SHSP_G_R_Q_R, `LD1SHSP_G_R_Q_F);
      if(!TE) (posedge G => (QN -: D)) = (`LD1SHSP_G_R_QN_R, `LD1SHSP_G_R_QN_F);
      if(TE) (posedge G => (QN -: TI)) = (`LD1SHSP_G_R_QN_R, `LD1SHSP_G_R_QN_F);
      if(!D && TI) (posedge G => (QN -: TE)) = (`LD1SHSP_G_R_QN_R, `LD1SHSP_G_R_QN_F);
      if(!TI && D) (posedge G => (QN +: TE)) = (`LD1SHSP_G_R_QN_R, `LD1SHSP_G_R_QN_F);

	$setuphold(negedge G &&& XorDTI_, posedge TE, `LD1SHSP_TE_G_SETUP_posedge_negedge, `LD1SHSP_TE_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& XorDTI_, negedge TE, `LD1SHSP_TE_G_SETUP_negedge_negedge, `LD1SHSP_TE_G_HOLD_negedge_negedge, Notifier);

	$setuphold(negedge G &&& TE, posedge TI, `LD1SHSP_TI_G_SETUP_posedge_negedge, `LD1SHSP_TI_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& TE, negedge TI, `LD1SHSP_TI_G_SETUP_negedge_negedge, `LD1SHSP_TI_G_HOLD_negedge_negedge, Notifier);

	$setuphold(negedge G &&& TEX, posedge D, `LD1SHSP_D_G_SETUP_posedge_negedge, `LD1SHSP_D_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& TEX, negedge D, `LD1SHSP_D_G_SETUP_negedge_negedge, `LD1SHSP_D_G_HOLD_negedge_negedge, Notifier);

      $width(posedge G, `LD1SHSP_G_PWH, 0, Notifier);
`else

     if (!D && G && TI) (TE -=> QN) = (`LD1SHSP_TE_F_QN_R,`LD1SHSP_TE_R_QN_F);
     if (D && G && !TI) (TE +=> QN) = (`LD1SHSP_TE_R_QN_R,`LD1SHSP_TE_F_QN_F);
      (TI -=> QN) = (`LD1SHSP_TI_F_QN_R,`LD1SHSP_TI_R_QN_F);
      (D -=> QN) = (`LD1SHSP_D_F_QN_R,`LD1SHSP_D_R_QN_F);
     if (!D && G && TI) (TE +=> Q) = (`LD1SHSP_TE_R_Q_R,`LD1SHSP_TE_F_Q_F);
      if (D && G && !TI) (TE -=> Q) = (`LD1SHSP_TE_F_Q_R,`LD1SHSP_TE_R_Q_F);
      (TI +=> Q) = (`LD1SHSP_TI_R_Q_R,`LD1SHSP_TI_F_Q_F);
      (D +=> Q) = (`LD1SHSP_D_R_Q_R,`LD1SHSP_D_F_Q_F);
      (posedge G => (Q +: Mux21DTITE_)) = (`LD1SHSP_G_R_Q_R, `LD1SHSP_G_R_Q_F);
      (posedge G => (QN -: Mux21DTITE_)) = (`LD1SHSP_G_R_QN_R, `LD1SHSP_G_R_QN_F);
 
        $setuphold(negedge G &&& XorDTI_, posedge TE, `LD1SHSP_TE_G_SETUP_posedge_negedge, `LD1SHSP_TE_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& XorDTI_, negedge TE, `LD1SHSP_TE_G_SETUP_negedge_negedge, `LD1SHSP_TE_G_HOLD_negedge_negedge, Notifier);
 
        $setuphold(negedge G &&& TE, posedge TI, `LD1SHSP_TI_G_SETUP_posedge_negedge, `LD1SHSP_TI_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& TE, negedge TI, `LD1SHSP_TI_G_SETUP_negedge_negedge, `LD1SHSP_TI_G_HOLD_negedge_negedge, Notifier);
 
        $setuphold(negedge G &&& TEX, posedge D, `LD1SHSP_D_G_SETUP_posedge_negedge, `LD1SHSP_D_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& TEX, negedge D, `LD1SHSP_D_G_SETUP_negedge_negedge, `LD1SHSP_D_G_HOLD_negedge_negedge, Notifier);
 
      $width(posedge G, `LD1SHSP_G_PWH, 0, Notifier);
`endif
   endspecify
`endif


endmodule // LD1SHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:45 and Version :1.1 //
 
//  START 
// CELL LD1SQHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD1SQHS_TE_F_Q_F 0.1
`define LD1SQHS_TE_R_Q_R 0.1
`define LD1SQHS_TE_F_Q_R 0.1
`define LD1SQHS_TE_R_Q_F 0.1
`define LD1SQHS_TI_F_Q_F 0.1
`define LD1SQHS_TI_R_Q_R 0.1
`define LD1SQHS_G_R_Q_R 0.1
`define LD1SQHS_G_R_Q_F 0.1
`define LD1SQHS_D_F_Q_F 0.1
`define LD1SQHS_D_R_Q_R 0.1
`define LD1SQHS_TE_G_HOLD_posedge_negedge 0.1
`define LD1SQHS_TE_G_HOLD_negedge_negedge 0.1
`define LD1SQHS_TE_G_SETUP_posedge_negedge 0.1
`define LD1SQHS_TE_G_SETUP_negedge_negedge 0.1
`define LD1SQHS_TI_G_HOLD_posedge_negedge 0.1
`define LD1SQHS_TI_G_HOLD_negedge_negedge 0.1
`define LD1SQHS_TI_G_SETUP_posedge_negedge 0.1
`define LD1SQHS_TI_G_SETUP_negedge_negedge 0.1
`define LD1SQHS_D_G_HOLD_posedge_negedge 0.1
`define LD1SQHS_D_G_HOLD_negedge_negedge 0.1
`define LD1SQHS_D_G_SETUP_posedge_negedge 0.1
`define LD1SQHS_D_G_SETUP_negedge_negedge 0.1
`define LD1SQHS_G_PWH 0.1

module LD1SQHS (Q, D, G, TI, TE);

   output Q;
   input D;
   input G;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_LD_P_NOTI u1 (IQ, Mux21DTITE_, G, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault

      if (!D && G && TI) (TE +=> Q) = (`LD1SQHS_TE_R_Q_R,`LD1SQHS_TE_F_Q_F);
      if (D && G && !TI) (TE -=> Q) = (`LD1SQHS_TE_F_Q_R,`LD1SQHS_TE_R_Q_F);
      if (G && TE) (TI +=> Q) = (`LD1SQHS_TI_R_Q_R,`LD1SQHS_TI_F_Q_F);
      if (G && !TE) (D +=> Q) = (`LD1SQHS_D_R_Q_R,`LD1SQHS_D_F_Q_F);
      if(!TE) (posedge G => (Q +: D)) = (`LD1SQHS_G_R_Q_R, `LD1SQHS_G_R_Q_F);
      if(TE) (posedge G => (Q +: TI)) = (`LD1SQHS_G_R_Q_R, `LD1SQHS_G_R_Q_F);
      if(!D && TI) (posedge G => (Q +: TE)) = (`LD1SQHS_G_R_Q_R, `LD1SQHS_G_R_Q_F);
      if(!TI && D) (posedge G => (Q -: TE)) = (`LD1SQHS_G_R_Q_R, `LD1SQHS_G_R_Q_F);

	$setuphold(negedge G &&& XorDTI_, posedge TE, `LD1SQHS_TE_G_SETUP_posedge_negedge, `LD1SQHS_TE_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& XorDTI_, negedge TE, `LD1SQHS_TE_G_SETUP_negedge_negedge, `LD1SQHS_TE_G_HOLD_negedge_negedge, Notifier);

	$setuphold(negedge G &&& TE, posedge TI, `LD1SQHS_TI_G_SETUP_posedge_negedge, `LD1SQHS_TI_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& TE, negedge TI, `LD1SQHS_TI_G_SETUP_negedge_negedge, `LD1SQHS_TI_G_HOLD_negedge_negedge, Notifier);

	$setuphold(negedge G &&& TEX, posedge D, `LD1SQHS_D_G_SETUP_posedge_negedge, `LD1SQHS_D_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& TEX, negedge D, `LD1SQHS_D_G_SETUP_negedge_negedge, `LD1SQHS_D_G_HOLD_negedge_negedge, Notifier);

      $width(posedge G, `LD1SQHS_G_PWH, 0, Notifier);
`else

     if (!D && G && TI) (TE +=> Q) = (`LD1SQHS_TE_R_Q_R,`LD1SQHS_TE_F_Q_F);
     if (D && G && !TI) (TE -=> Q) = (`LD1SQHS_TE_F_Q_R,`LD1SQHS_TE_R_Q_F);
      (TI +=> Q) = (`LD1SQHS_TI_R_Q_R,`LD1SQHS_TI_F_Q_F);
      (D +=> Q) = (`LD1SQHS_D_R_Q_R,`LD1SQHS_D_F_Q_F);
      (posedge G => (Q +: Mux21DTITE_)) = (`LD1SQHS_G_R_Q_R, `LD1SQHS_G_R_Q_F);
 
        $setuphold(negedge G &&& XorDTI_, posedge TE, `LD1SQHS_TE_G_SETUP_posedge_negedge, `LD1SQHS_TE_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& XorDTI_, negedge TE, `LD1SQHS_TE_G_SETUP_negedge_negedge, `LD1SQHS_TE_G_HOLD_negedge_negedge, Notifier);
 
        $setuphold(negedge G &&& TE, posedge TI, `LD1SQHS_TI_G_SETUP_posedge_negedge, `LD1SQHS_TI_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& TE, negedge TI, `LD1SQHS_TI_G_SETUP_negedge_negedge, `LD1SQHS_TI_G_HOLD_negedge_negedge, Notifier);
 
        $setuphold(negedge G &&& TEX, posedge D, `LD1SQHS_D_G_SETUP_posedge_negedge, `LD1SQHS_D_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& TEX, negedge D, `LD1SQHS_D_G_SETUP_negedge_negedge, `LD1SQHS_D_G_HOLD_negedge_negedge, Notifier);
 
      $width(posedge G, `LD1SQHS_G_PWH, 0, Notifier);
`endif
   endspecify
`endif


endmodule // LD1SQHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:45 and Version :1.1 //
 
//  START 
// CELL LD1SQHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD1SQHSP_TE_F_Q_F 0.1
`define LD1SQHSP_TE_R_Q_R 0.1
`define LD1SQHSP_TE_F_Q_R 0.1
`define LD1SQHSP_TE_R_Q_F 0.1
`define LD1SQHSP_TI_F_Q_F 0.1
`define LD1SQHSP_TI_R_Q_R 0.1
`define LD1SQHSP_G_R_Q_R 0.1
`define LD1SQHSP_G_R_Q_F 0.1
`define LD1SQHSP_D_F_Q_F 0.1
`define LD1SQHSP_D_R_Q_R 0.1
`define LD1SQHSP_TE_G_HOLD_posedge_negedge 0.1
`define LD1SQHSP_TE_G_HOLD_negedge_negedge 0.1
`define LD1SQHSP_TE_G_SETUP_posedge_negedge 0.1
`define LD1SQHSP_TE_G_SETUP_negedge_negedge 0.1
`define LD1SQHSP_TI_G_HOLD_posedge_negedge 0.1
`define LD1SQHSP_TI_G_HOLD_negedge_negedge 0.1
`define LD1SQHSP_TI_G_SETUP_posedge_negedge 0.1
`define LD1SQHSP_TI_G_SETUP_negedge_negedge 0.1
`define LD1SQHSP_D_G_HOLD_posedge_negedge 0.1
`define LD1SQHSP_D_G_HOLD_negedge_negedge 0.1
`define LD1SQHSP_D_G_SETUP_posedge_negedge 0.1
`define LD1SQHSP_D_G_SETUP_negedge_negedge 0.1
`define LD1SQHSP_G_PWH 0.1

module LD1SQHSP (Q, D, G, TI, TE);

   output Q;
   input D;
   input G;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_LD_P_NOTI u1 (IQ, Mux21DTITE_, G, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault

      if (!D && G && TI) (TE +=> Q) = (`LD1SQHSP_TE_R_Q_R,`LD1SQHSP_TE_F_Q_F);
      if (D && G && !TI) (TE -=> Q) = (`LD1SQHSP_TE_F_Q_R,`LD1SQHSP_TE_R_Q_F);
      if (G && TE) (TI +=> Q) = (`LD1SQHSP_TI_R_Q_R,`LD1SQHSP_TI_F_Q_F);
      if (G && !TE) (D +=> Q) = (`LD1SQHSP_D_R_Q_R,`LD1SQHSP_D_F_Q_F);
      if(!TE) (posedge G => (Q +: D)) = (`LD1SQHSP_G_R_Q_R, `LD1SQHSP_G_R_Q_F);
      if(TE) (posedge G => (Q +: TI)) = (`LD1SQHSP_G_R_Q_R, `LD1SQHSP_G_R_Q_F);
      if(!D && TI) (posedge G => (Q +: TE)) = (`LD1SQHSP_G_R_Q_R, `LD1SQHSP_G_R_Q_F);
      if(!TI && D) (posedge G => (Q -: TE)) = (`LD1SQHSP_G_R_Q_R, `LD1SQHSP_G_R_Q_F);

	$setuphold(negedge G &&& XorDTI_, posedge TE, `LD1SQHSP_TE_G_SETUP_posedge_negedge, `LD1SQHSP_TE_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& XorDTI_, negedge TE, `LD1SQHSP_TE_G_SETUP_negedge_negedge, `LD1SQHSP_TE_G_HOLD_negedge_negedge, Notifier);

	$setuphold(negedge G &&& TE, posedge TI, `LD1SQHSP_TI_G_SETUP_posedge_negedge, `LD1SQHSP_TI_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& TE, negedge TI, `LD1SQHSP_TI_G_SETUP_negedge_negedge, `LD1SQHSP_TI_G_HOLD_negedge_negedge, Notifier);

	$setuphold(negedge G &&& TEX, posedge D, `LD1SQHSP_D_G_SETUP_posedge_negedge, `LD1SQHSP_D_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& TEX, negedge D, `LD1SQHSP_D_G_SETUP_negedge_negedge, `LD1SQHSP_D_G_HOLD_negedge_negedge, Notifier);

      $width(posedge G, `LD1SQHSP_G_PWH, 0, Notifier);
`else

     if (!D && G && TI) (TE +=> Q) = (`LD1SQHSP_TE_R_Q_R,`LD1SQHSP_TE_F_Q_F);
     if (D && G && !TI) (TE -=> Q) = (`LD1SQHSP_TE_F_Q_R,`LD1SQHSP_TE_R_Q_F);
      (TI +=> Q) = (`LD1SQHSP_TI_R_Q_R,`LD1SQHSP_TI_F_Q_F);
      (D +=> Q) = (`LD1SQHSP_D_R_Q_R,`LD1SQHSP_D_F_Q_F);
      (posedge G => (Q +: Mux21DTITE_)) = (`LD1SQHSP_G_R_Q_R, `LD1SQHSP_G_R_Q_F);
 
        $setuphold(negedge G &&& XorDTI_, posedge TE, `LD1SQHSP_TE_G_SETUP_posedge_negedge, `LD1SQHSP_TE_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& XorDTI_, negedge TE, `LD1SQHSP_TE_G_SETUP_negedge_negedge, `LD1SQHSP_TE_G_HOLD_negedge_negedge, Notifier);
 
        $setuphold(negedge G &&& TE, posedge TI, `LD1SQHSP_TI_G_SETUP_posedge_negedge, `LD1SQHSP_TI_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& TE, negedge TI, `LD1SQHSP_TI_G_SETUP_negedge_negedge, `LD1SQHSP_TI_G_HOLD_negedge_negedge, Notifier);
 
        $setuphold(negedge G &&& TEX, posedge D, `LD1SQHSP_D_G_SETUP_posedge_negedge, `LD1SQHSP_D_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& TEX, negedge D, `LD1SQHSP_D_G_SETUP_negedge_negedge, `LD1SQHSP_D_G_HOLD_negedge_negedge, Notifier);
 
      $width(posedge G, `LD1SQHSP_G_PWH, 0, Notifier);
`endif
   endspecify
`endif


endmodule // LD1SQHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:45 and Version :1.1 //
 
//  START 
// CELL LD1SQHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD1SQHSX4_TE_F_Q_F 0.1
`define LD1SQHSX4_TE_R_Q_R 0.1
`define LD1SQHSX4_TE_F_Q_R 0.1
`define LD1SQHSX4_TE_R_Q_F 0.1
`define LD1SQHSX4_TI_F_Q_F 0.1
`define LD1SQHSX4_TI_R_Q_R 0.1
`define LD1SQHSX4_G_R_Q_R 0.1
`define LD1SQHSX4_G_R_Q_F 0.1
`define LD1SQHSX4_D_F_Q_F 0.1
`define LD1SQHSX4_D_R_Q_R 0.1
`define LD1SQHSX4_TE_G_HOLD_posedge_negedge 0.1
`define LD1SQHSX4_TE_G_HOLD_negedge_negedge 0.1
`define LD1SQHSX4_TE_G_SETUP_posedge_negedge 0.1
`define LD1SQHSX4_TE_G_SETUP_negedge_negedge 0.1
`define LD1SQHSX4_TI_G_HOLD_posedge_negedge 0.1
`define LD1SQHSX4_TI_G_HOLD_negedge_negedge 0.1
`define LD1SQHSX4_TI_G_SETUP_posedge_negedge 0.1
`define LD1SQHSX4_TI_G_SETUP_negedge_negedge 0.1
`define LD1SQHSX4_D_G_HOLD_posedge_negedge 0.1
`define LD1SQHSX4_D_G_HOLD_negedge_negedge 0.1
`define LD1SQHSX4_D_G_SETUP_posedge_negedge 0.1
`define LD1SQHSX4_D_G_SETUP_negedge_negedge 0.1
`define LD1SQHSX4_G_PWH 0.1

module LD1SQHSX4 (Q, D, G, TI, TE);

   output Q;
   input D;
   input G;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_LD_P_NOTI u1 (IQ, Mux21DTITE_, G, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault

      if (!D && G && TI) (TE +=> Q) = (`LD1SQHSX4_TE_R_Q_R,`LD1SQHSX4_TE_F_Q_F);
      if (D && G && !TI) (TE -=> Q) = (`LD1SQHSX4_TE_F_Q_R,`LD1SQHSX4_TE_R_Q_F);
      if (G && TE) (TI +=> Q) = (`LD1SQHSX4_TI_R_Q_R,`LD1SQHSX4_TI_F_Q_F);
      if (G && !TE) (D +=> Q) = (`LD1SQHSX4_D_R_Q_R,`LD1SQHSX4_D_F_Q_F);
      if(!TE) (posedge G => (Q +: D)) = (`LD1SQHSX4_G_R_Q_R, `LD1SQHSX4_G_R_Q_F);
      if(TE) (posedge G => (Q +: TI)) = (`LD1SQHSX4_G_R_Q_R, `LD1SQHSX4_G_R_Q_F);
      if(!D && TI) (posedge G => (Q +: TE)) = (`LD1SQHSX4_G_R_Q_R, `LD1SQHSX4_G_R_Q_F);
      if(!TI && D) (posedge G => (Q -: TE)) = (`LD1SQHSX4_G_R_Q_R, `LD1SQHSX4_G_R_Q_F);

	$setuphold(negedge G &&& XorDTI_, posedge TE, `LD1SQHSX4_TE_G_SETUP_posedge_negedge, `LD1SQHSX4_TE_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& XorDTI_, negedge TE, `LD1SQHSX4_TE_G_SETUP_negedge_negedge, `LD1SQHSX4_TE_G_HOLD_negedge_negedge, Notifier);

	$setuphold(negedge G &&& TE, posedge TI, `LD1SQHSX4_TI_G_SETUP_posedge_negedge, `LD1SQHSX4_TI_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& TE, negedge TI, `LD1SQHSX4_TI_G_SETUP_negedge_negedge, `LD1SQHSX4_TI_G_HOLD_negedge_negedge, Notifier);

	$setuphold(negedge G &&& TEX, posedge D, `LD1SQHSX4_D_G_SETUP_posedge_negedge, `LD1SQHSX4_D_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& TEX, negedge D, `LD1SQHSX4_D_G_SETUP_negedge_negedge, `LD1SQHSX4_D_G_HOLD_negedge_negedge, Notifier);

      $width(posedge G, `LD1SQHSX4_G_PWH, 0, Notifier);
`else

     if (!D && G && TI) (TE +=> Q) = (`LD1SQHSX4_TE_R_Q_R,`LD1SQHSX4_TE_F_Q_F);
     if (D && G && !TI) (TE -=> Q) = (`LD1SQHSX4_TE_F_Q_R,`LD1SQHSX4_TE_R_Q_F);
      (TI +=> Q) = (`LD1SQHSX4_TI_R_Q_R,`LD1SQHSX4_TI_F_Q_F);
      (D +=> Q) = (`LD1SQHSX4_D_R_Q_R,`LD1SQHSX4_D_F_Q_F);
      (posedge G => (Q +: Mux21DTITE_)) = (`LD1SQHSX4_G_R_Q_R, `LD1SQHSX4_G_R_Q_F);
 
        $setuphold(negedge G &&& XorDTI_, posedge TE, `LD1SQHSX4_TE_G_SETUP_posedge_negedge, `LD1SQHSX4_TE_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& XorDTI_, negedge TE, `LD1SQHSX4_TE_G_SETUP_negedge_negedge, `LD1SQHSX4_TE_G_HOLD_negedge_negedge, Notifier);
 
        $setuphold(negedge G &&& TE, posedge TI, `LD1SQHSX4_TI_G_SETUP_posedge_negedge, `LD1SQHSX4_TI_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& TE, negedge TI, `LD1SQHSX4_TI_G_SETUP_negedge_negedge, `LD1SQHSX4_TI_G_HOLD_negedge_negedge, Notifier);
 
        $setuphold(negedge G &&& TEX, posedge D, `LD1SQHSX4_D_G_SETUP_posedge_negedge, `LD1SQHSX4_D_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& TEX, negedge D, `LD1SQHSX4_D_G_SETUP_negedge_negedge, `LD1SQHSX4_D_G_HOLD_negedge_negedge, Notifier);
 
      $width(posedge G, `LD1SQHSX4_G_PWH, 0, Notifier);
`endif
   endspecify
`endif


endmodule // LD1SQHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:45 and Version :1.1 //
 
//  START 
// CELL LD2HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD2HS_GN_F_QN_F 0.1
`define LD2HS_GN_F_QN_R 0.1
`define LD2HS_D_F_QN_R 0.1
`define LD2HS_D_R_QN_F 0.1
`define LD2HS_GN_F_Q_R 0.1
`define LD2HS_GN_F_Q_F 0.1
`define LD2HS_D_F_Q_F 0.1
`define LD2HS_D_R_Q_R 0.1
`define LD2HS_GN_PWL 0.1
`define LD2HS_D_GN_SETUP_posedge_posedge 0.1
`define LD2HS_D_GN_SETUP_negedge_posedge 0.1
`define LD2HS_D_GN_HOLD_posedge_posedge 0.1
`define LD2HS_D_GN_HOLD_negedge_posedge 0.1

module LD2HS (Q, QN, D, GN);

   output Q;
   output QN;
   input D;
   input GN;


   reg Notifier;


   U_LD_N_NOTI u0 (   // Verilog Seq UDP
      IQ, D, GN, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   specify

      if (!GN) (D -=> QN) = (`LD2HS_D_F_QN_R,`LD2HS_D_R_QN_F);
      if (!GN) (D +=> Q) = (`LD2HS_D_R_Q_R,`LD2HS_D_F_Q_F);
      (negedge GN => (Q +: D)) = (`LD2HS_GN_F_Q_R, `LD2HS_GN_F_Q_F);
      (negedge GN => (QN -: D)) = (`LD2HS_GN_F_QN_R, `LD2HS_GN_F_QN_F);

	$setuphold(posedge GN, posedge D, `LD2HS_D_GN_SETUP_posedge_posedge, `LD2HS_D_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN, negedge D, `LD2HS_D_GN_SETUP_negedge_posedge, `LD2HS_D_GN_HOLD_negedge_posedge, Notifier);

      $width(negedge GN, `LD2HS_GN_PWL, 0, Notifier);

   endspecify
`endif


endmodule // LD2HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:49 and Version :1.1 //
 
//  START 
// CELL LD2HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD2HSP_GN_F_QN_F 0.1
`define LD2HSP_GN_F_QN_R 0.1
`define LD2HSP_D_F_QN_R 0.1
`define LD2HSP_D_R_QN_F 0.1
`define LD2HSP_GN_F_Q_R 0.1
`define LD2HSP_GN_F_Q_F 0.1
`define LD2HSP_D_F_Q_F 0.1
`define LD2HSP_D_R_Q_R 0.1
`define LD2HSP_GN_PWL 0.1
`define LD2HSP_D_GN_SETUP_posedge_posedge 0.1
`define LD2HSP_D_GN_SETUP_negedge_posedge 0.1
`define LD2HSP_D_GN_HOLD_posedge_posedge 0.1
`define LD2HSP_D_GN_HOLD_negedge_posedge 0.1

module LD2HSP (Q, QN, D, GN);

   output Q;
   output QN;
   input D;
   input GN;


   reg Notifier;


   U_LD_N_NOTI u0 (   // Verilog Seq UDP
      IQ, D, GN, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   specify

      if (!GN) (D -=> QN) = (`LD2HSP_D_F_QN_R,`LD2HSP_D_R_QN_F);
      if (!GN) (D +=> Q) = (`LD2HSP_D_R_Q_R,`LD2HSP_D_F_Q_F);
      (negedge GN => (Q +: D)) = (`LD2HSP_GN_F_Q_R, `LD2HSP_GN_F_Q_F);
      (negedge GN => (QN -: D)) = (`LD2HSP_GN_F_QN_R, `LD2HSP_GN_F_QN_F);

	$setuphold(posedge GN, posedge D, `LD2HSP_D_GN_SETUP_posedge_posedge, `LD2HSP_D_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN, negedge D, `LD2HSP_D_GN_SETUP_negedge_posedge, `LD2HSP_D_GN_HOLD_negedge_posedge, Notifier);

      $width(negedge GN, `LD2HSP_GN_PWL, 0, Notifier);

   endspecify
`endif


endmodule // LD2HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:49 and Version :1.1 //
 
//  START 
// CELL LD2QHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD2QHS_GN_F_Q_R 0.1
`define LD2QHS_GN_F_Q_F 0.1
`define LD2QHS_D_F_Q_F 0.1
`define LD2QHS_D_R_Q_R 0.1
`define LD2QHS_D_GN_HOLD_posedge_posedge 0.1
`define LD2QHS_D_GN_HOLD_negedge_posedge 0.1
`define LD2QHS_D_GN_SETUP_posedge_posedge 0.1
`define LD2QHS_D_GN_SETUP_negedge_posedge 0.1
`define LD2QHS_GN_PWL 0.1

module LD2QHS (Q, D, GN);

   output Q;
   input D;
   input GN;


   reg Notifier;


   U_LD_N_NOTI u0 (IQ, D, GN, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify

      if (!GN) (D +=> Q) = (`LD2QHS_D_R_Q_R,`LD2QHS_D_F_Q_F);
      (negedge GN => (Q +: D)) = (`LD2QHS_GN_F_Q_R, `LD2QHS_GN_F_Q_F);

	$setuphold(posedge GN, posedge D, `LD2QHS_D_GN_SETUP_posedge_posedge, `LD2QHS_D_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN, negedge D, `LD2QHS_D_GN_SETUP_negedge_posedge, `LD2QHS_D_GN_HOLD_negedge_posedge, Notifier);

      $width(negedge GN, `LD2QHS_GN_PWL, 0, Notifier);

   endspecify
`endif


endmodule // LD2QHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:51 and Version :1.1 //
 
//  START 
// CELL LD2QHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD2QHSP_GN_F_Q_R 0.1
`define LD2QHSP_GN_F_Q_F 0.1
`define LD2QHSP_D_F_Q_F 0.1
`define LD2QHSP_D_R_Q_R 0.1
`define LD2QHSP_D_GN_HOLD_posedge_posedge 0.1
`define LD2QHSP_D_GN_HOLD_negedge_posedge 0.1
`define LD2QHSP_D_GN_SETUP_posedge_posedge 0.1
`define LD2QHSP_D_GN_SETUP_negedge_posedge 0.1
`define LD2QHSP_GN_PWL 0.1

module LD2QHSP (Q, D, GN);

   output Q;
   input D;
   input GN;


   reg Notifier;


   U_LD_N_NOTI u0 (IQ, D, GN, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify

      if (!GN) (D +=> Q) = (`LD2QHSP_D_R_Q_R,`LD2QHSP_D_F_Q_F);
      (negedge GN => (Q +: D)) = (`LD2QHSP_GN_F_Q_R, `LD2QHSP_GN_F_Q_F);

	$setuphold(posedge GN, posedge D, `LD2QHSP_D_GN_SETUP_posedge_posedge, `LD2QHSP_D_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN, negedge D, `LD2QHSP_D_GN_SETUP_negedge_posedge, `LD2QHSP_D_GN_HOLD_negedge_posedge, Notifier);

      $width(negedge GN, `LD2QHSP_GN_PWL, 0, Notifier);

   endspecify
`endif


endmodule // LD2QHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:51 and Version :1.1 //
 
//  START 
// CELL LD2QHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD2QHSX4_GN_F_Q_R 0.1
`define LD2QHSX4_GN_F_Q_F 0.1
`define LD2QHSX4_D_F_Q_F 0.1
`define LD2QHSX4_D_R_Q_R 0.1
`define LD2QHSX4_D_GN_HOLD_posedge_posedge 0.1
`define LD2QHSX4_D_GN_HOLD_negedge_posedge 0.1
`define LD2QHSX4_D_GN_SETUP_posedge_posedge 0.1
`define LD2QHSX4_D_GN_SETUP_negedge_posedge 0.1
`define LD2QHSX4_GN_PWL 0.1

module LD2QHSX4 (Q, D, GN);

   output Q;
   input D;
   input GN;


   reg Notifier;


   U_LD_N_NOTI u0 (IQ, D, GN, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify

      if (!GN) (D +=> Q) = (`LD2QHSX4_D_R_Q_R,`LD2QHSX4_D_F_Q_F);
      (negedge GN => (Q +: D)) = (`LD2QHSX4_GN_F_Q_R, `LD2QHSX4_GN_F_Q_F);

	$setuphold(posedge GN, posedge D, `LD2QHSX4_D_GN_SETUP_posedge_posedge, `LD2QHSX4_D_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN, negedge D, `LD2QHSX4_D_GN_SETUP_negedge_posedge, `LD2QHSX4_D_GN_HOLD_negedge_posedge, Notifier);

      $width(negedge GN, `LD2QHSX4_GN_PWL, 0, Notifier);

   endspecify
`endif


endmodule // LD2QHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:51 and Version :1.1 //
 
//  START 
// CELL LD2SHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD2SHS_TE_F_QN_R 0.1
`define LD2SHS_TE_R_QN_F 0.1
`define LD2SHS_TE_F_QN_F 0.1
`define LD2SHS_TE_R_QN_R 0.1
`define LD2SHS_TI_F_QN_R 0.1
`define LD2SHS_TI_R_QN_F 0.1
`define LD2SHS_GN_F_QN_F 0.1
`define LD2SHS_GN_F_QN_R 0.1
`define LD2SHS_D_F_QN_R 0.1
`define LD2SHS_D_R_QN_F 0.1
`define LD2SHS_TE_F_Q_F 0.1
`define LD2SHS_TE_R_Q_R 0.1
`define LD2SHS_TE_F_Q_R 0.1
`define LD2SHS_TE_R_Q_F 0.1
`define LD2SHS_TI_F_Q_F 0.1
`define LD2SHS_TI_R_Q_R 0.1
`define LD2SHS_GN_F_Q_R 0.1
`define LD2SHS_GN_F_Q_F 0.1
`define LD2SHS_D_F_Q_F 0.1
`define LD2SHS_D_R_Q_R 0.1
`define LD2SHS_GN_PWL 0.1
`define LD2SHS_D_GN_SETUP_posedge_posedge 0.1
`define LD2SHS_D_GN_SETUP_negedge_posedge 0.1
`define LD2SHS_D_GN_HOLD_posedge_posedge 0.1
`define LD2SHS_D_GN_HOLD_negedge_posedge 0.1
`define LD2SHS_TI_GN_SETUP_posedge_posedge 0.1
`define LD2SHS_TI_GN_SETUP_negedge_posedge 0.1
`define LD2SHS_TI_GN_HOLD_posedge_posedge 0.1
`define LD2SHS_TI_GN_HOLD_negedge_posedge 0.1
`define LD2SHS_TE_GN_SETUP_posedge_posedge 0.1
`define LD2SHS_TE_GN_SETUP_negedge_posedge 0.1
`define LD2SHS_TE_GN_HOLD_posedge_posedge 0.1
`define LD2SHS_TE_GN_HOLD_negedge_posedge 0.1

module LD2SHS (Q, QN, D, GN, TI, TE);

   output Q;
   output QN;
   input D;
   input GN;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_LD_N_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, GN, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault

      if (!D && !GN && TI) (TE -=> QN) = (`LD2SHS_TE_F_QN_R,`LD2SHS_TE_R_QN_F);
      if (D && !GN && !TI) (TE +=> QN) = (`LD2SHS_TE_R_QN_R,`LD2SHS_TE_F_QN_F);
      if (!GN && TE) (TI -=> QN) = (`LD2SHS_TI_F_QN_R,`LD2SHS_TI_R_QN_F);
      if (!GN && !TE) (D -=> QN) = (`LD2SHS_D_F_QN_R,`LD2SHS_D_R_QN_F);
      if (!D && !GN && TI) (TE +=> Q) = (`LD2SHS_TE_R_Q_R,`LD2SHS_TE_F_Q_F);
      if (D && !GN && !TI) (TE -=> Q) = (`LD2SHS_TE_F_Q_R,`LD2SHS_TE_R_Q_F);
      if (!GN && TE) (TI +=> Q) = (`LD2SHS_TI_R_Q_R,`LD2SHS_TI_F_Q_F);
      if (!GN && !TE) (D +=> Q) = (`LD2SHS_D_R_Q_R,`LD2SHS_D_F_Q_F);
      if(!TE) (negedge GN => (Q +: D)) = (`LD2SHS_GN_F_Q_R, `LD2SHS_GN_F_Q_F);
      if(TE) (negedge GN => (Q +: TI)) = (`LD2SHS_GN_F_Q_R, `LD2SHS_GN_F_Q_F);
      if(!D && TI) (negedge GN => (Q +: TE)) = (`LD2SHS_GN_F_Q_R, `LD2SHS_GN_F_Q_F);
      if(!TI && D) (negedge GN => (Q -: TE)) = (`LD2SHS_GN_F_Q_R, `LD2SHS_GN_F_Q_F);
      if(!TE) (negedge GN => (QN -: D)) = (`LD2SHS_GN_F_QN_R, `LD2SHS_GN_F_QN_F);
      if(TE) (negedge GN => (QN -: TI)) = (`LD2SHS_GN_F_QN_R, `LD2SHS_GN_F_QN_F);
      if(!D && TI) (negedge GN => (QN -: TE)) = (`LD2SHS_GN_F_QN_R, `LD2SHS_GN_F_QN_F);
      if(!TI && D) (negedge GN => (QN +: TE)) = (`LD2SHS_GN_F_QN_R, `LD2SHS_GN_F_QN_F);

	$setuphold(posedge GN &&& XorDTI_, posedge TE, `LD2SHS_TE_GN_SETUP_posedge_posedge, `LD2SHS_TE_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& XorDTI_, negedge TE, `LD2SHS_TE_GN_SETUP_negedge_posedge, `LD2SHS_TE_GN_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge GN &&& TE, posedge TI, `LD2SHS_TI_GN_SETUP_posedge_posedge, `LD2SHS_TI_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& TE, negedge TI, `LD2SHS_TI_GN_SETUP_negedge_posedge, `LD2SHS_TI_GN_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge GN &&& TEX, posedge D, `LD2SHS_D_GN_SETUP_posedge_posedge, `LD2SHS_D_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& TEX, negedge D, `LD2SHS_D_GN_SETUP_negedge_posedge, `LD2SHS_D_GN_HOLD_negedge_posedge, Notifier);

      $width(negedge GN, `LD2SHS_GN_PWL, 0, Notifier);
`else

     if (!D && !GN && TI) (TE -=> QN) = (`LD2SHS_TE_F_QN_R,`LD2SHS_TE_R_QN_F);
     if (D && !GN && !TI) (TE +=> QN) = (`LD2SHS_TE_R_QN_R,`LD2SHS_TE_F_QN_F);
      (TI -=> QN) = (`LD2SHS_TI_F_QN_R,`LD2SHS_TI_R_QN_F);
      (D -=> QN) = (`LD2SHS_D_F_QN_R,`LD2SHS_D_R_QN_F);
     if (!D && !GN && TI) (TE +=> Q) = (`LD2SHS_TE_R_Q_R,`LD2SHS_TE_F_Q_F);
      if (D && !GN && !TI) (TE -=> Q) = (`LD2SHS_TE_F_Q_R,`LD2SHS_TE_R_Q_F);
      (TI +=> Q) = (`LD2SHS_TI_R_Q_R,`LD2SHS_TI_F_Q_F);
      (D +=> Q) = (`LD2SHS_D_R_Q_R,`LD2SHS_D_F_Q_F);
      (negedge GN => (Q +: Mux21DTITE_)) = (`LD2SHS_GN_F_Q_R, `LD2SHS_GN_F_Q_F);
      (negedge GN => (QN -: Mux21DTITE_)) = (`LD2SHS_GN_F_QN_R, `LD2SHS_GN_F_QN_F);
 
        $setuphold(posedge GN &&& XorDTI_, posedge TE, `LD2SHS_TE_GN_SETUP_posedge_posedge, `LD2SHS_TE_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& XorDTI_, negedge TE, `LD2SHS_TE_GN_SETUP_negedge_posedge, `LD2SHS_TE_GN_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge GN &&& TE, posedge TI, `LD2SHS_TI_GN_SETUP_posedge_posedge, `LD2SHS_TI_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& TE, negedge TI, `LD2SHS_TI_GN_SETUP_negedge_posedge, `LD2SHS_TI_GN_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge GN &&& TEX, posedge D, `LD2SHS_D_GN_SETUP_posedge_posedge, `LD2SHS_D_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& TEX, negedge D, `LD2SHS_D_GN_SETUP_negedge_posedge, `LD2SHS_D_GN_HOLD_negedge_posedge, Notifier);
 
      $width(negedge GN, `LD2SHS_GN_PWL, 0, Notifier);
`endif
   endspecify
`endif


endmodule // LD2SHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:57 and Version :1.1 //
 
//  START 
// CELL LD2SQHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD2SQHS_TE_F_Q_F 0.1
`define LD2SQHS_TE_R_Q_R 0.1
`define LD2SQHS_TE_F_Q_R 0.1
`define LD2SQHS_TE_R_Q_F 0.1
`define LD2SQHS_TI_F_Q_F 0.1
`define LD2SQHS_TI_R_Q_R 0.1
`define LD2SQHS_GN_F_Q_R 0.1
`define LD2SQHS_GN_F_Q_F 0.1
`define LD2SQHS_D_F_Q_F 0.1
`define LD2SQHS_D_R_Q_R 0.1
`define LD2SQHS_TE_GN_HOLD_posedge_posedge 0.1
`define LD2SQHS_TE_GN_HOLD_negedge_posedge 0.1
`define LD2SQHS_TE_GN_SETUP_posedge_posedge 0.1
`define LD2SQHS_TE_GN_SETUP_negedge_posedge 0.1
`define LD2SQHS_TI_GN_HOLD_posedge_posedge 0.1
`define LD2SQHS_TI_GN_HOLD_negedge_posedge 0.1
`define LD2SQHS_TI_GN_SETUP_posedge_posedge 0.1
`define LD2SQHS_TI_GN_SETUP_negedge_posedge 0.1
`define LD2SQHS_D_GN_HOLD_posedge_posedge 0.1
`define LD2SQHS_D_GN_HOLD_negedge_posedge 0.1
`define LD2SQHS_D_GN_SETUP_posedge_posedge 0.1
`define LD2SQHS_D_GN_SETUP_negedge_posedge 0.1
`define LD2SQHS_GN_PWL 0.1

module LD2SQHS (Q, D, GN, TI, TE);

   output Q;
   input D;
   input GN;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_LD_N_NOTI u1 (IQ, Mux21DTITE_, GN, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault

      if (!D && !GN && TI) (TE +=> Q) = (`LD2SQHS_TE_R_Q_R,`LD2SQHS_TE_F_Q_F);
      if (D && !GN && !TI) (TE -=> Q) = (`LD2SQHS_TE_F_Q_R,`LD2SQHS_TE_R_Q_F);
      if (!GN && TE) (TI +=> Q) = (`LD2SQHS_TI_R_Q_R,`LD2SQHS_TI_F_Q_F);
      if (!GN && !TE) (D +=> Q) = (`LD2SQHS_D_R_Q_R,`LD2SQHS_D_F_Q_F);
      if(!TE) (negedge GN => (Q +: D)) = (`LD2SQHS_GN_F_Q_R, `LD2SQHS_GN_F_Q_F);
      if(TE) (negedge GN => (Q +: TI)) = (`LD2SQHS_GN_F_Q_R, `LD2SQHS_GN_F_Q_F);
      if(!D && TI) (negedge GN => (Q +: TE)) = (`LD2SQHS_GN_F_Q_R, `LD2SQHS_GN_F_Q_F);
      if(!TI && D) (negedge GN => (Q -: TE)) = (`LD2SQHS_GN_F_Q_R, `LD2SQHS_GN_F_Q_F);

	$setuphold(posedge GN &&& XorDTI_, posedge TE, `LD2SQHS_TE_GN_SETUP_posedge_posedge, `LD2SQHS_TE_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& XorDTI_, negedge TE, `LD2SQHS_TE_GN_SETUP_negedge_posedge, `LD2SQHS_TE_GN_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge GN &&& TE, posedge TI, `LD2SQHS_TI_GN_SETUP_posedge_posedge, `LD2SQHS_TI_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& TE, negedge TI, `LD2SQHS_TI_GN_SETUP_negedge_posedge, `LD2SQHS_TI_GN_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge GN &&& TEX, posedge D, `LD2SQHS_D_GN_SETUP_posedge_posedge, `LD2SQHS_D_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& TEX, negedge D, `LD2SQHS_D_GN_SETUP_negedge_posedge, `LD2SQHS_D_GN_HOLD_negedge_posedge, Notifier);

      $width(negedge GN, `LD2SQHS_GN_PWL, 0, Notifier);
`else

     if (!D && !GN && TI) (TE +=> Q) = (`LD2SQHS_TE_R_Q_R,`LD2SQHS_TE_F_Q_F);
      if (D && !GN && !TI) (TE -=> Q) = (`LD2SQHS_TE_F_Q_R,`LD2SQHS_TE_R_Q_F);
      (TI +=> Q) = (`LD2SQHS_TI_R_Q_R,`LD2SQHS_TI_F_Q_F);
      (D +=> Q) = (`LD2SQHS_D_R_Q_R,`LD2SQHS_D_F_Q_F);
      (negedge GN => (Q +: Mux21DTITE_)) = (`LD2SQHS_GN_F_Q_R, `LD2SQHS_GN_F_Q_F);
 
        $setuphold(posedge GN &&& XorDTI_, posedge TE, `LD2SQHS_TE_GN_SETUP_posedge_posedge, `LD2SQHS_TE_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& XorDTI_, negedge TE, `LD2SQHS_TE_GN_SETUP_negedge_posedge, `LD2SQHS_TE_GN_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge GN &&& TE, posedge TI, `LD2SQHS_TI_GN_SETUP_posedge_posedge, `LD2SQHS_TI_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& TE, negedge TI, `LD2SQHS_TI_GN_SETUP_negedge_posedge, `LD2SQHS_TI_GN_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge GN &&& TEX, posedge D, `LD2SQHS_D_GN_SETUP_posedge_posedge, `LD2SQHS_D_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& TEX, negedge D, `LD2SQHS_D_GN_SETUP_negedge_posedge, `LD2SQHS_D_GN_HOLD_negedge_posedge, Notifier);
 
      $width(negedge GN, `LD2SQHS_GN_PWL, 0, Notifier);
`endif
   endspecify
`endif


endmodule // LD2SQHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:57 and Version :1.1 //
 
//  START 
// CELL LD2SQHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD2SQHSP_TE_F_Q_F 0.1
`define LD2SQHSP_TE_R_Q_R 0.1
`define LD2SQHSP_TE_F_Q_R 0.1
`define LD2SQHSP_TE_R_Q_F 0.1
`define LD2SQHSP_TI_F_Q_F 0.1
`define LD2SQHSP_TI_R_Q_R 0.1
`define LD2SQHSP_GN_F_Q_R 0.1
`define LD2SQHSP_GN_F_Q_F 0.1
`define LD2SQHSP_D_F_Q_F 0.1
`define LD2SQHSP_D_R_Q_R 0.1
`define LD2SQHSP_TE_GN_HOLD_posedge_posedge 0.1
`define LD2SQHSP_TE_GN_HOLD_negedge_posedge 0.1
`define LD2SQHSP_TE_GN_SETUP_posedge_posedge 0.1
`define LD2SQHSP_TE_GN_SETUP_negedge_posedge 0.1
`define LD2SQHSP_TI_GN_HOLD_posedge_posedge 0.1
`define LD2SQHSP_TI_GN_HOLD_negedge_posedge 0.1
`define LD2SQHSP_TI_GN_SETUP_posedge_posedge 0.1
`define LD2SQHSP_TI_GN_SETUP_negedge_posedge 0.1
`define LD2SQHSP_D_GN_HOLD_posedge_posedge 0.1
`define LD2SQHSP_D_GN_HOLD_negedge_posedge 0.1
`define LD2SQHSP_D_GN_SETUP_posedge_posedge 0.1
`define LD2SQHSP_D_GN_SETUP_negedge_posedge 0.1
`define LD2SQHSP_GN_PWL 0.1

module LD2SQHSP (Q, D, GN, TI, TE);

   output Q;
   input D;
   input GN;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_LD_N_NOTI u1 (IQ, Mux21DTITE_, GN, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault

      if (!D && !GN && TI) (TE +=> Q) = (`LD2SQHSP_TE_R_Q_R,`LD2SQHSP_TE_F_Q_F);
      if (D && !GN && !TI) (TE -=> Q) = (`LD2SQHSP_TE_F_Q_R,`LD2SQHSP_TE_R_Q_F);
      if (!GN && TE) (TI +=> Q) = (`LD2SQHSP_TI_R_Q_R,`LD2SQHSP_TI_F_Q_F);
      if (!GN && !TE) (D +=> Q) = (`LD2SQHSP_D_R_Q_R,`LD2SQHSP_D_F_Q_F);
      if(!TE) (negedge GN => (Q +: D)) = (`LD2SQHSP_GN_F_Q_R, `LD2SQHSP_GN_F_Q_F);
      if(TE) (negedge GN => (Q +: TI)) = (`LD2SQHSP_GN_F_Q_R, `LD2SQHSP_GN_F_Q_F);
      if(!D && TI) (negedge GN => (Q +: TE)) = (`LD2SQHSP_GN_F_Q_R, `LD2SQHSP_GN_F_Q_F);
      if(!TI && D) (negedge GN => (Q -: TE)) = (`LD2SQHSP_GN_F_Q_R, `LD2SQHSP_GN_F_Q_F);

	$setuphold(posedge GN &&& XorDTI_, posedge TE, `LD2SQHSP_TE_GN_SETUP_posedge_posedge, `LD2SQHSP_TE_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& XorDTI_, negedge TE, `LD2SQHSP_TE_GN_SETUP_negedge_posedge, `LD2SQHSP_TE_GN_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge GN &&& TE, posedge TI, `LD2SQHSP_TI_GN_SETUP_posedge_posedge, `LD2SQHSP_TI_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& TE, negedge TI, `LD2SQHSP_TI_GN_SETUP_negedge_posedge, `LD2SQHSP_TI_GN_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge GN &&& TEX, posedge D, `LD2SQHSP_D_GN_SETUP_posedge_posedge, `LD2SQHSP_D_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& TEX, negedge D, `LD2SQHSP_D_GN_SETUP_negedge_posedge, `LD2SQHSP_D_GN_HOLD_negedge_posedge, Notifier);

      $width(negedge GN, `LD2SQHSP_GN_PWL, 0, Notifier);
`else

     if (!D && !GN && TI) (TE +=> Q) = (`LD2SQHSP_TE_R_Q_R,`LD2SQHSP_TE_F_Q_F);
      if (D && !GN && !TI) (TE -=> Q) = (`LD2SQHSP_TE_F_Q_R,`LD2SQHSP_TE_R_Q_F);
      (TI +=> Q) = (`LD2SQHSP_TI_R_Q_R,`LD2SQHSP_TI_F_Q_F);
      (D +=> Q) = (`LD2SQHSP_D_R_Q_R,`LD2SQHSP_D_F_Q_F);
      (negedge GN => (Q +: Mux21DTITE_)) = (`LD2SQHSP_GN_F_Q_R, `LD2SQHSP_GN_F_Q_F);
 
        $setuphold(posedge GN &&& XorDTI_, posedge TE, `LD2SQHSP_TE_GN_SETUP_posedge_posedge, `LD2SQHSP_TE_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& XorDTI_, negedge TE, `LD2SQHSP_TE_GN_SETUP_negedge_posedge, `LD2SQHSP_TE_GN_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge GN &&& TE, posedge TI, `LD2SQHSP_TI_GN_SETUP_posedge_posedge, `LD2SQHSP_TI_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& TE, negedge TI, `LD2SQHSP_TI_GN_SETUP_negedge_posedge, `LD2SQHSP_TI_GN_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge GN &&& TEX, posedge D, `LD2SQHSP_D_GN_SETUP_posedge_posedge, `LD2SQHSP_D_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& TEX, negedge D, `LD2SQHSP_D_GN_SETUP_negedge_posedge, `LD2SQHSP_D_GN_HOLD_negedge_posedge, Notifier);
 
      $width(negedge GN, `LD2SQHSP_GN_PWL, 0, Notifier);
`endif
   endspecify
`endif


endmodule // LD2SQHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:57 and Version :1.1 //
 
//  START 
// CELL LD2SQHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD2SQHSX4_TE_F_Q_F 0.1
`define LD2SQHSX4_TE_R_Q_R 0.1
`define LD2SQHSX4_TE_F_Q_R 0.1
`define LD2SQHSX4_TE_R_Q_F 0.1
`define LD2SQHSX4_TI_F_Q_F 0.1
`define LD2SQHSX4_TI_R_Q_R 0.1
`define LD2SQHSX4_GN_F_Q_R 0.1
`define LD2SQHSX4_GN_F_Q_F 0.1
`define LD2SQHSX4_D_F_Q_F 0.1
`define LD2SQHSX4_D_R_Q_R 0.1
`define LD2SQHSX4_TE_GN_HOLD_posedge_posedge 0.1
`define LD2SQHSX4_TE_GN_HOLD_negedge_posedge 0.1
`define LD2SQHSX4_TE_GN_SETUP_posedge_posedge 0.1
`define LD2SQHSX4_TE_GN_SETUP_negedge_posedge 0.1
`define LD2SQHSX4_TI_GN_HOLD_posedge_posedge 0.1
`define LD2SQHSX4_TI_GN_HOLD_negedge_posedge 0.1
`define LD2SQHSX4_TI_GN_SETUP_posedge_posedge 0.1
`define LD2SQHSX4_TI_GN_SETUP_negedge_posedge 0.1
`define LD2SQHSX4_D_GN_HOLD_posedge_posedge 0.1
`define LD2SQHSX4_D_GN_HOLD_negedge_posedge 0.1
`define LD2SQHSX4_D_GN_SETUP_posedge_posedge 0.1
`define LD2SQHSX4_D_GN_SETUP_negedge_posedge 0.1
`define LD2SQHSX4_GN_PWL 0.1

module LD2SQHSX4 (Q, D, GN, TI, TE);

   output Q;
   input D;
   input GN;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_LD_N_NOTI u1 (IQ, Mux21DTITE_, GN, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   xor  (XorDTI_, D, TI);
   specify
`ifdef verifault

      if (!D && !GN && TI) (TE +=> Q) = (`LD2SQHSX4_TE_R_Q_R,`LD2SQHSX4_TE_F_Q_F);
      if (D && !GN && !TI) (TE -=> Q) = (`LD2SQHSX4_TE_F_Q_R,`LD2SQHSX4_TE_R_Q_F);
      if (!GN && TE) (TI +=> Q) = (`LD2SQHSX4_TI_R_Q_R,`LD2SQHSX4_TI_F_Q_F);
      if (!GN && !TE) (D +=> Q) = (`LD2SQHSX4_D_R_Q_R,`LD2SQHSX4_D_F_Q_F);
      if(!TE) (negedge GN => (Q +: D)) = (`LD2SQHSX4_GN_F_Q_R, `LD2SQHSX4_GN_F_Q_F);
      if(TE) (negedge GN => (Q +: TI)) = (`LD2SQHSX4_GN_F_Q_R, `LD2SQHSX4_GN_F_Q_F);
      if(!D && TI) (negedge GN => (Q +: TE)) = (`LD2SQHSX4_GN_F_Q_R, `LD2SQHSX4_GN_F_Q_F);
      if(!TI && D) (negedge GN => (Q -: TE)) = (`LD2SQHSX4_GN_F_Q_R, `LD2SQHSX4_GN_F_Q_F);

	$setuphold(posedge GN &&& XorDTI_, posedge TE, `LD2SQHSX4_TE_GN_SETUP_posedge_posedge, `LD2SQHSX4_TE_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& XorDTI_, negedge TE, `LD2SQHSX4_TE_GN_SETUP_negedge_posedge, `LD2SQHSX4_TE_GN_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge GN &&& TE, posedge TI, `LD2SQHSX4_TI_GN_SETUP_posedge_posedge, `LD2SQHSX4_TI_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& TE, negedge TI, `LD2SQHSX4_TI_GN_SETUP_negedge_posedge, `LD2SQHSX4_TI_GN_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge GN &&& TEX, posedge D, `LD2SQHSX4_D_GN_SETUP_posedge_posedge, `LD2SQHSX4_D_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& TEX, negedge D, `LD2SQHSX4_D_GN_SETUP_negedge_posedge, `LD2SQHSX4_D_GN_HOLD_negedge_posedge, Notifier);

      $width(negedge GN, `LD2SQHSX4_GN_PWL, 0, Notifier);
`else

     if (!D && !GN && TI) (TE +=> Q) = (`LD2SQHSX4_TE_R_Q_R,`LD2SQHSX4_TE_F_Q_F);
      if (D && !GN && !TI) (TE -=> Q) = (`LD2SQHSX4_TE_F_Q_R,`LD2SQHSX4_TE_R_Q_F);
      (TI +=> Q) = (`LD2SQHSX4_TI_R_Q_R,`LD2SQHSX4_TI_F_Q_F);
      (D +=> Q) = (`LD2SQHSX4_D_R_Q_R,`LD2SQHSX4_D_F_Q_F);
      (negedge GN => (Q +: Mux21DTITE_)) = (`LD2SQHSX4_GN_F_Q_R, `LD2SQHSX4_GN_F_Q_F);
 
        $setuphold(posedge GN &&& XorDTI_, posedge TE, `LD2SQHSX4_TE_GN_SETUP_posedge_posedge, `LD2SQHSX4_TE_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& XorDTI_, negedge TE, `LD2SQHSX4_TE_GN_SETUP_negedge_posedge, `LD2SQHSX4_TE_GN_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge GN &&& TE, posedge TI, `LD2SQHSX4_TI_GN_SETUP_posedge_posedge, `LD2SQHSX4_TI_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& TE, negedge TI, `LD2SQHSX4_TI_GN_SETUP_negedge_posedge, `LD2SQHSX4_TI_GN_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge GN &&& TEX, posedge D, `LD2SQHSX4_D_GN_SETUP_posedge_posedge, `LD2SQHSX4_D_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& TEX, negedge D, `LD2SQHSX4_D_GN_SETUP_negedge_posedge, `LD2SQHSX4_D_GN_HOLD_negedge_posedge, Notifier);
 
      $width(negedge GN, `LD2SQHSX4_GN_PWL, 0, Notifier);
`endif
   endspecify
`endif


endmodule // LD2SQHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:17:57 and Version :1.1 //
 
//  START 
// CELL LD3HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD3HS_CD_F_QN_R 0.1
`define LD3HS_CD_R_QN_F 0.1
`define LD3HS_G_R_QN_F 0.1
`define LD3HS_G_R_QN_R 0.1
`define LD3HS_D_F_QN_R 0.1
`define LD3HS_D_R_QN_F 0.1
`define LD3HS_CD_F_Q_F 0.1
`define LD3HS_CD_R_Q_R 0.1
`define LD3HS_G_R_Q_R 0.1
`define LD3HS_G_R_Q_F 0.1
`define LD3HS_D_F_Q_F 0.1
`define LD3HS_D_R_Q_R 0.1
`define LD3HS_CD_G_REM_posedge_negedge 0.1
`define LD3HS_CD_G_REC_posedge_negedge 0.1
`define LD3HS_CD_PWL 0.1
`define LD3HS_G_PWH 0.1
`define LD3HS_D_G_SETUP_posedge_negedge 0.1
`define LD3HS_D_G_SETUP_negedge_negedge 0.1
`define LD3HS_D_G_HOLD_posedge_negedge 0.1
`define LD3HS_D_G_HOLD_negedge_negedge 0.1

module LD3HS (Q, QN, D, G, CD);

   output Q;
   output QN;
   input D;
   input G;
   input CD;


   reg Notifier;


   U_LD_P_RN_NOTI u0 (   // Verilog Seq UDP
      IQ,  D, G, CD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   not  (GX, G);
   specify
`ifdef verifault

      if (G && CD) (D -=> QN) = (`LD3HS_D_F_QN_R,`LD3HS_D_R_QN_F);
      if (G && CD) (D +=> Q) = (`LD3HS_D_R_Q_R,`LD3HS_D_F_Q_F);
      (posedge G => (Q +: D)) = (`LD3HS_G_R_Q_R, `LD3HS_G_R_Q_F);
      (posedge G => (QN -: D)) = (`LD3HS_G_R_QN_R, `LD3HS_G_R_QN_F);
      if(D && G) (posedge CD => (Q +: 1'b1)) = (`LD3HS_CD_R_Q_R,`LD3HS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD3HS_CD_R_Q_R,`LD3HS_CD_F_Q_F);
      if(D && G) (posedge CD => (QN +: 1'b0)) = (`LD3HS_CD_F_QN_R,`LD3HS_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`LD3HS_CD_F_QN_R,`LD3HS_CD_R_QN_F);

	$setuphold(negedge G &&& CD, posedge D, `LD3HS_D_G_SETUP_posedge_negedge, `LD3HS_D_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& CD, negedge D, `LD3HS_D_G_SETUP_negedge_negedge, `LD3HS_D_G_HOLD_negedge_negedge, Notifier);

      $width(posedge G, `LD3HS_G_PWH, 0, Notifier);
      $width(negedge CD, `LD3HS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, negedge G &&& D, `LD3HS_CD_G_REC_posedge_negedge, Notifier);

	$hold(negedge G &&& D, posedge CD, `LD3HS_CD_G_REM_posedge_negedge, Notifier);

`else

      (D -=> QN) = (`LD3HS_D_F_QN_R,`LD3HS_D_R_QN_F);
      (D +=> Q) = (`LD3HS_D_R_Q_R,`LD3HS_D_F_Q_F);
      (posedge G => (Q +: D)) = (`LD3HS_G_R_Q_R, `LD3HS_G_R_Q_F);
      (posedge G => (QN -: D)) = (`LD3HS_G_R_QN_R, `LD3HS_G_R_QN_F);
      (posedge CD => (Q +: 1'b1)) = (`LD3HS_CD_R_Q_R,`LD3HS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD3HS_CD_R_Q_R,`LD3HS_CD_F_Q_F);
      (posedge CD => (QN +: 1'b0)) = (`LD3HS_CD_F_QN_R,`LD3HS_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`LD3HS_CD_F_QN_R,`LD3HS_CD_R_QN_F);
 
        $setuphold(negedge G &&& CD, posedge D, `LD3HS_D_G_SETUP_posedge_negedge, `LD3HS_D_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& CD, negedge D, `LD3HS_D_G_SETUP_negedge_negedge, `LD3HS_D_G_HOLD_negedge_negedge, Notifier);
 
      $width(posedge G, `LD3HS_G_PWH, 0, Notifier);
      $width(negedge CD, `LD3HS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, negedge G &&& D, `LD3HS_CD_G_REC_posedge_negedge, Notifier);
 
        $hold(negedge G &&& D, posedge CD, `LD3HS_CD_G_REM_posedge_negedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD3HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:01 and Version :1.1 //
 
//  START 
// CELL LD3HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD3HSP_CD_F_QN_R 0.1
`define LD3HSP_CD_R_QN_F 0.1
`define LD3HSP_G_R_QN_F 0.1
`define LD3HSP_G_R_QN_R 0.1
`define LD3HSP_D_F_QN_R 0.1
`define LD3HSP_D_R_QN_F 0.1
`define LD3HSP_CD_F_Q_F 0.1
`define LD3HSP_CD_R_Q_R 0.1
`define LD3HSP_G_R_Q_R 0.1
`define LD3HSP_G_R_Q_F 0.1
`define LD3HSP_D_F_Q_F 0.1
`define LD3HSP_D_R_Q_R 0.1
`define LD3HSP_CD_G_REM_posedge_negedge 0.1
`define LD3HSP_CD_G_REC_posedge_negedge 0.1
`define LD3HSP_CD_PWL 0.1
`define LD3HSP_G_PWH 0.1
`define LD3HSP_D_G_SETUP_posedge_negedge 0.1
`define LD3HSP_D_G_SETUP_negedge_negedge 0.1
`define LD3HSP_D_G_HOLD_posedge_negedge 0.1
`define LD3HSP_D_G_HOLD_negedge_negedge 0.1

module LD3HSP (Q, QN, D, G, CD);

   output Q;
   output QN;
   input D;
   input G;
   input CD;


   reg Notifier;


   U_LD_P_RN_NOTI u0 (   // Verilog Seq UDP
      IQ,  D, G, CD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   not  (GX, G);
   specify
`ifdef verifault

      if (G && CD) (D -=> QN) = (`LD3HSP_D_F_QN_R,`LD3HSP_D_R_QN_F);
      if (G && CD) (D +=> Q) = (`LD3HSP_D_R_Q_R,`LD3HSP_D_F_Q_F);
      (posedge G => (Q +: D)) = (`LD3HSP_G_R_Q_R, `LD3HSP_G_R_Q_F);
      (posedge G => (QN -: D)) = (`LD3HSP_G_R_QN_R, `LD3HSP_G_R_QN_F);
      if(D && G) (posedge CD => (Q +: 1'b1)) = (`LD3HSP_CD_R_Q_R,`LD3HSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD3HSP_CD_R_Q_R,`LD3HSP_CD_F_Q_F);
      if(D && G) (posedge CD => (QN +: 1'b0)) = (`LD3HSP_CD_F_QN_R,`LD3HSP_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`LD3HSP_CD_F_QN_R,`LD3HSP_CD_R_QN_F);

	$setuphold(negedge G &&& CD, posedge D, `LD3HSP_D_G_SETUP_posedge_negedge, `LD3HSP_D_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& CD, negedge D, `LD3HSP_D_G_SETUP_negedge_negedge, `LD3HSP_D_G_HOLD_negedge_negedge, Notifier);

      $width(posedge G, `LD3HSP_G_PWH, 0, Notifier);
      $width(negedge CD, `LD3HSP_CD_PWL, 0, Notifier);
	$recovery(posedge CD, negedge G &&& D, `LD3HSP_CD_G_REC_posedge_negedge, Notifier);

	$hold(negedge G &&& D, posedge CD, `LD3HSP_CD_G_REM_posedge_negedge, Notifier);

`else

      (D -=> QN) = (`LD3HSP_D_F_QN_R,`LD3HSP_D_R_QN_F);
      (D +=> Q) = (`LD3HSP_D_R_Q_R,`LD3HSP_D_F_Q_F);
      (posedge G => (Q +: D)) = (`LD3HSP_G_R_Q_R, `LD3HSP_G_R_Q_F);
      (posedge G => (QN -: D)) = (`LD3HSP_G_R_QN_R, `LD3HSP_G_R_QN_F);
      (posedge CD => (Q +: 1'b1)) = (`LD3HSP_CD_R_Q_R,`LD3HSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD3HSP_CD_R_Q_R,`LD3HSP_CD_F_Q_F);
      (posedge CD => (QN +: 1'b0)) = (`LD3HSP_CD_F_QN_R,`LD3HSP_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`LD3HSP_CD_F_QN_R,`LD3HSP_CD_R_QN_F);
 
        $setuphold(negedge G &&& CD, posedge D, `LD3HSP_D_G_SETUP_posedge_negedge, `LD3HSP_D_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& CD, negedge D, `LD3HSP_D_G_SETUP_negedge_negedge, `LD3HSP_D_G_HOLD_negedge_negedge, Notifier);
 
      $width(posedge G, `LD3HSP_G_PWH, 0, Notifier);
      $width(negedge CD, `LD3HSP_CD_PWL, 0, Notifier);
        $recovery(posedge CD, negedge G &&& D, `LD3HSP_CD_G_REC_posedge_negedge, Notifier);
 
        $hold(negedge G &&& D, posedge CD, `LD3HSP_CD_G_REM_posedge_negedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD3HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:01 and Version :1.1 //
 
//  START 
// CELL LD3QHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD3QHS_CD_F_Q_F 0.1
`define LD3QHS_CD_R_Q_R 0.1
`define LD3QHS_G_R_Q_R 0.1
`define LD3QHS_G_R_Q_F 0.1
`define LD3QHS_D_F_Q_F 0.1
`define LD3QHS_D_R_Q_R 0.1
`define LD3QHS_D_G_HOLD_posedge_negedge 0.1
`define LD3QHS_D_G_HOLD_negedge_negedge 0.1
`define LD3QHS_D_G_SETUP_posedge_negedge 0.1
`define LD3QHS_D_G_SETUP_negedge_negedge 0.1
`define LD3QHS_G_PWH 0.1
`define LD3QHS_CD_PWL 0.1
`define LD3QHS_CD_G_REC_posedge_negedge 0.1
`define LD3QHS_CD_G_REM_posedge_negedge 0.1

module LD3QHS (Q, D, G, CD);

   output Q;
   input D;
   input G;
   input CD;


   reg Notifier;


   U_LD_P_RN_NOTI u0 (IQ, D, G, CD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   not  (GX, G);
   specify
`ifdef verifault

      if (G && CD) (D +=> Q) = (`LD3QHS_D_R_Q_R,`LD3QHS_D_F_Q_F);
      if(CD) (posedge G => (Q +: D)) = (`LD3QHS_G_R_Q_R, `LD3QHS_G_R_Q_F);
      if(D && G) (posedge CD => (Q +: 1'b1)) = (`LD3QHS_CD_R_Q_R,`LD3QHS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD3QHS_CD_R_Q_R,`LD3QHS_CD_F_Q_F);

	$setuphold(negedge G &&& CD, posedge D, `LD3QHS_D_G_SETUP_posedge_negedge, `LD3QHS_D_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& CD, negedge D, `LD3QHS_D_G_SETUP_negedge_negedge, `LD3QHS_D_G_HOLD_negedge_negedge, Notifier);

      $width(posedge G, `LD3QHS_G_PWH, 0, Notifier);
      $width(negedge CD, `LD3QHS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, negedge G &&& D, `LD3QHS_CD_G_REC_posedge_negedge, Notifier);

	$hold(negedge G &&& D, posedge CD, `LD3QHS_CD_G_REM_posedge_negedge, Notifier);

`else

      (D +=> Q) = (`LD3QHS_D_R_Q_R,`LD3QHS_D_F_Q_F);
      (posedge G => (Q +: D)) = (`LD3QHS_G_R_Q_R, `LD3QHS_G_R_Q_F);
      (posedge CD => (Q +: 1'b1)) = (`LD3QHS_CD_R_Q_R,`LD3QHS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD3QHS_CD_R_Q_R,`LD3QHS_CD_F_Q_F);
 
        $setuphold(negedge G &&& CD, posedge D, `LD3QHS_D_G_SETUP_posedge_negedge, `LD3QHS_D_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& CD, negedge D, `LD3QHS_D_G_SETUP_negedge_negedge, `LD3QHS_D_G_HOLD_negedge_negedge, Notifier);
 
      $width(posedge G, `LD3QHS_G_PWH, 0, Notifier);
      $width(negedge CD, `LD3QHS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, negedge G &&& D, `LD3QHS_CD_G_REC_posedge_negedge, Notifier);
 
        $hold(negedge G &&& D, posedge CD, `LD3QHS_CD_G_REM_posedge_negedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD3QHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:03 and Version :1.1 //
 
//  START 
// CELL LD3QHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD3QHSP_CD_F_Q_F 0.1
`define LD3QHSP_CD_R_Q_R 0.1
`define LD3QHSP_G_R_Q_R 0.1
`define LD3QHSP_G_R_Q_F 0.1
`define LD3QHSP_D_F_Q_F 0.1
`define LD3QHSP_D_R_Q_R 0.1
`define LD3QHSP_D_G_HOLD_posedge_negedge 0.1
`define LD3QHSP_D_G_HOLD_negedge_negedge 0.1
`define LD3QHSP_D_G_SETUP_posedge_negedge 0.1
`define LD3QHSP_D_G_SETUP_negedge_negedge 0.1
`define LD3QHSP_G_PWH 0.1
`define LD3QHSP_CD_PWL 0.1
`define LD3QHSP_CD_G_REC_posedge_negedge 0.1
`define LD3QHSP_CD_G_REM_posedge_negedge 0.1

module LD3QHSP (Q, D, G, CD);

   output Q;
   input D;
   input G;
   input CD;


   reg Notifier;


   U_LD_P_RN_NOTI u0 (IQ, D, G, CD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   not  (GX, G);
   specify
`ifdef verifault

      if (G && CD) (D +=> Q) = (`LD3QHSP_D_R_Q_R,`LD3QHSP_D_F_Q_F);
      if(CD) (posedge G => (Q +: D)) = (`LD3QHSP_G_R_Q_R, `LD3QHSP_G_R_Q_F);
      if(D && G) (posedge CD => (Q +: 1'b1)) = (`LD3QHSP_CD_R_Q_R,`LD3QHSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD3QHSP_CD_R_Q_R,`LD3QHSP_CD_F_Q_F);

	$setuphold(negedge G &&& CD, posedge D, `LD3QHSP_D_G_SETUP_posedge_negedge, `LD3QHSP_D_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& CD, negedge D, `LD3QHSP_D_G_SETUP_negedge_negedge, `LD3QHSP_D_G_HOLD_negedge_negedge, Notifier);

      $width(posedge G, `LD3QHSP_G_PWH, 0, Notifier);
      $width(negedge CD, `LD3QHSP_CD_PWL, 0, Notifier);
	$recovery(posedge CD, negedge G &&& D, `LD3QHSP_CD_G_REC_posedge_negedge, Notifier);

	$hold(negedge G &&& D, posedge CD, `LD3QHSP_CD_G_REM_posedge_negedge, Notifier);

`else

      (D +=> Q) = (`LD3QHSP_D_R_Q_R,`LD3QHSP_D_F_Q_F);
      (posedge G => (Q +: D)) = (`LD3QHSP_G_R_Q_R, `LD3QHSP_G_R_Q_F);
      (posedge CD => (Q +: 1'b1)) = (`LD3QHSP_CD_R_Q_R,`LD3QHSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD3QHSP_CD_R_Q_R,`LD3QHSP_CD_F_Q_F);
 
        $setuphold(negedge G &&& CD, posedge D, `LD3QHSP_D_G_SETUP_posedge_negedge, `LD3QHSP_D_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& CD, negedge D, `LD3QHSP_D_G_SETUP_negedge_negedge, `LD3QHSP_D_G_HOLD_negedge_negedge, Notifier);
 
      $width(posedge G, `LD3QHSP_G_PWH, 0, Notifier);
      $width(negedge CD, `LD3QHSP_CD_PWL, 0, Notifier);
        $recovery(posedge CD, negedge G &&& D, `LD3QHSP_CD_G_REC_posedge_negedge, Notifier);
 
        $hold(negedge G &&& D, posedge CD, `LD3QHSP_CD_G_REM_posedge_negedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD3QHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:03 and Version :1.1 //
 
//  START 
// CELL LD3QHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD3QHSX4_CD_F_Q_F 0.1
`define LD3QHSX4_CD_R_Q_R 0.1
`define LD3QHSX4_G_R_Q_R 0.1
`define LD3QHSX4_G_R_Q_F 0.1
`define LD3QHSX4_D_F_Q_F 0.1
`define LD3QHSX4_D_R_Q_R 0.1
`define LD3QHSX4_D_G_HOLD_posedge_negedge 0.1
`define LD3QHSX4_D_G_HOLD_negedge_negedge 0.1
`define LD3QHSX4_D_G_SETUP_posedge_negedge 0.1
`define LD3QHSX4_D_G_SETUP_negedge_negedge 0.1
`define LD3QHSX4_G_PWH 0.1
`define LD3QHSX4_CD_PWL 0.1
`define LD3QHSX4_CD_G_REC_posedge_negedge 0.1
`define LD3QHSX4_CD_G_REM_posedge_negedge 0.1

module LD3QHSX4 (Q, D, G, CD);

   output Q;
   input D;
   input G;
   input CD;


   reg Notifier;


   U_LD_P_RN_NOTI u0 (IQ, D, G, CD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   not  (GX, G);
   specify
`ifdef verifault

      if (G && CD) (D +=> Q) = (`LD3QHSX4_D_R_Q_R,`LD3QHSX4_D_F_Q_F);
      if(CD) (posedge G => (Q +: D)) = (`LD3QHSX4_G_R_Q_R, `LD3QHSX4_G_R_Q_F);
      if(D && G) (posedge CD => (Q +: 1'b1)) = (`LD3QHSX4_CD_R_Q_R,`LD3QHSX4_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD3QHSX4_CD_R_Q_R,`LD3QHSX4_CD_F_Q_F);

	$setuphold(negedge G &&& CD, posedge D, `LD3QHSX4_D_G_SETUP_posedge_negedge, `LD3QHSX4_D_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& CD, negedge D, `LD3QHSX4_D_G_SETUP_negedge_negedge, `LD3QHSX4_D_G_HOLD_negedge_negedge, Notifier);

      $width(posedge G, `LD3QHSX4_G_PWH, 0, Notifier);
      $width(negedge CD, `LD3QHSX4_CD_PWL, 0, Notifier);
	$recovery(posedge CD, negedge G &&& D, `LD3QHSX4_CD_G_REC_posedge_negedge, Notifier);

	$hold(negedge G &&& D, posedge CD, `LD3QHSX4_CD_G_REM_posedge_negedge, Notifier);

`else

      (D +=> Q) = (`LD3QHSX4_D_R_Q_R,`LD3QHSX4_D_F_Q_F);
      (posedge G => (Q +: D)) = (`LD3QHSX4_G_R_Q_R, `LD3QHSX4_G_R_Q_F);
      (posedge CD => (Q +: 1'b1)) = (`LD3QHSX4_CD_R_Q_R,`LD3QHSX4_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD3QHSX4_CD_R_Q_R,`LD3QHSX4_CD_F_Q_F);
 
        $setuphold(negedge G &&& CD, posedge D, `LD3QHSX4_D_G_SETUP_posedge_negedge, `LD3QHSX4_D_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& CD, negedge D, `LD3QHSX4_D_G_SETUP_negedge_negedge, `LD3QHSX4_D_G_HOLD_negedge_negedge, Notifier);
 
      $width(posedge G, `LD3QHSX4_G_PWH, 0, Notifier);
      $width(negedge CD, `LD3QHSX4_CD_PWL, 0, Notifier);
        $recovery(posedge CD, negedge G &&& D, `LD3QHSX4_CD_G_REC_posedge_negedge, Notifier);
 
        $hold(negedge G &&& D, posedge CD, `LD3QHSX4_CD_G_REM_posedge_negedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD3QHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:03 and Version :1.1 //
 
//  START 
// CELL LD3SHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD3SHS_TE_F_QN_R 0.1
`define LD3SHS_TE_R_QN_F 0.1
`define LD3SHS_TE_F_QN_F 0.1
`define LD3SHS_TE_R_QN_R 0.1
`define LD3SHS_TI_F_QN_R 0.1
`define LD3SHS_TI_R_QN_F 0.1
`define LD3SHS_CD_F_QN_R 0.1
`define LD3SHS_CD_R_QN_F 0.1
`define LD3SHS_G_R_QN_F 0.1
`define LD3SHS_G_R_QN_R 0.1
`define LD3SHS_D_F_QN_R 0.1
`define LD3SHS_D_R_QN_F 0.1
`define LD3SHS_TE_F_Q_F 0.1
`define LD3SHS_TE_R_Q_R 0.1
`define LD3SHS_TE_F_Q_R 0.1
`define LD3SHS_TE_R_Q_F 0.1
`define LD3SHS_TI_F_Q_F 0.1
`define LD3SHS_TI_R_Q_R 0.1
`define LD3SHS_CD_F_Q_F 0.1
`define LD3SHS_CD_R_Q_R 0.1
`define LD3SHS_G_R_Q_R 0.1
`define LD3SHS_G_R_Q_F 0.1
`define LD3SHS_D_F_Q_F 0.1
`define LD3SHS_D_R_Q_R 0.1
`define LD3SHS_CD_G_REM_posedge_negedge 0.1
`define LD3SHS_CD_G_REC_posedge_negedge 0.1
`define LD3SHS_CD_PWL 0.1
`define LD3SHS_G_PWH 0.1
`define LD3SHS_D_G_SETUP_posedge_negedge 0.1
`define LD3SHS_D_G_SETUP_negedge_negedge 0.1
`define LD3SHS_D_G_HOLD_posedge_negedge 0.1
`define LD3SHS_D_G_HOLD_negedge_negedge 0.1
`define LD3SHS_TI_G_SETUP_posedge_negedge 0.1
`define LD3SHS_TI_G_SETUP_negedge_negedge 0.1
`define LD3SHS_TI_G_HOLD_posedge_negedge 0.1
`define LD3SHS_TI_G_HOLD_negedge_negedge 0.1
`define LD3SHS_TE_G_SETUP_posedge_negedge 0.1
`define LD3SHS_TE_G_SETUP_negedge_negedge 0.1
`define LD3SHS_TE_G_HOLD_posedge_negedge 0.1
`define LD3SHS_TE_G_HOLD_negedge_negedge 0.1

module LD3SHS (Q, QN, D, G, CD, TI, TE);

   output Q;
   output QN;
   input D;
   input G;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_LD_P_RN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, G, CD, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   not  (GX, G);
   not  (TEX, TE);
   and  (AndCDTEX_, CD, TEX);
   and  (AndCDTE_, CD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   specify
`ifdef verifault
      if (!D && G && TI) (TE -=> QN) = (`LD3SHS_TE_F_QN_R,`LD3SHS_TE_R_QN_F);
      if (D && G && !TI) (TE +=> QN) = (`LD3SHS_TE_R_QN_R,`LD3SHS_TE_F_QN_F);
      if (G && CD && TE) (TI -=> QN) = (`LD3SHS_TI_F_QN_R,`LD3SHS_TI_R_QN_F);
      if (G && CD && !TE) (D -=> QN) = (`LD3SHS_D_F_QN_R,`LD3SHS_D_R_QN_F);
      if (!D && G && TI) (TE +=> Q) = (`LD3SHS_TE_R_Q_R,`LD3SHS_TE_F_Q_F);
      if (D && G && !TI) (TE -=> Q) = (`LD3SHS_TE_F_Q_R,`LD3SHS_TE_R_Q_F);
      if (G && CD && TE) (TI +=> Q) = (`LD3SHS_TI_R_Q_R,`LD3SHS_TI_F_Q_F);
      if (G && CD && !TE) (D +=> Q) = (`LD3SHS_D_R_Q_R,`LD3SHS_D_F_Q_F);
      if(!TE) (posedge G => (Q +: D)) = (`LD3SHS_G_R_Q_R, `LD3SHS_G_R_Q_F);
      if(TE) (posedge G => (Q +: TI)) = (`LD3SHS_G_R_Q_R, `LD3SHS_G_R_Q_F);
      if(!D && TI) (posedge G => (Q +: TE)) = (`LD3SHS_G_R_Q_R, `LD3SHS_G_R_Q_F);
      if(!TI && D) (posedge G => (Q -: TE)) = (`LD3SHS_G_R_Q_R, `LD3SHS_G_R_Q_F);
      if(!TE) (posedge G => (QN -: D)) = (`LD3SHS_G_R_QN_R, `LD3SHS_G_R_QN_F);
      if(TE) (posedge G => (QN -: TI)) = (`LD3SHS_G_R_QN_R, `LD3SHS_G_R_QN_F);
      if(!D && TI) (posedge G => (QN -: TE)) = (`LD3SHS_G_R_QN_R, `LD3SHS_G_R_QN_F);
      if(!TI && D) (posedge G => (QN +: TE)) = (`LD3SHS_G_R_QN_R, `LD3SHS_G_R_QN_F);
      if(D && G && !TE || G && TI && TE) (posedge CD => (Q +: 1'b1)) = (`LD3SHS_CD_R_Q_R,`LD3SHS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD3SHS_CD_R_Q_R,`LD3SHS_CD_F_Q_F);
      if(D && G && !TE || G && TI && TE) (posedge CD => (QN +: 1'b0)) = (`LD3SHS_CD_F_QN_R,`LD3SHS_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`LD3SHS_CD_F_QN_R,`LD3SHS_CD_R_QN_F);

	$setuphold(negedge G &&& AndXorDTI_CD_, posedge TE, `LD3SHS_TE_G_SETUP_posedge_negedge, `LD3SHS_TE_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& AndXorDTI_CD_, negedge TE, `LD3SHS_TE_G_SETUP_negedge_negedge, `LD3SHS_TE_G_HOLD_negedge_negedge, Notifier);

	$setuphold(negedge G &&& AndCDTE_, posedge TI, `LD3SHS_TI_G_SETUP_posedge_negedge, `LD3SHS_TI_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& AndCDTE_, negedge TI, `LD3SHS_TI_G_SETUP_negedge_negedge, `LD3SHS_TI_G_HOLD_negedge_negedge, Notifier);

	$setuphold(negedge G &&& AndCDTEX_, posedge D, `LD3SHS_D_G_SETUP_posedge_negedge, `LD3SHS_D_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& AndCDTEX_, negedge D, `LD3SHS_D_G_SETUP_negedge_negedge, `LD3SHS_D_G_HOLD_negedge_negedge, Notifier);

      $width(posedge G, `LD3SHS_G_PWH, 0, Notifier);
      $width(negedge CD, `LD3SHS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, negedge G &&& Mux21DTITE_, `LD3SHS_CD_G_REC_posedge_negedge, Notifier);

	$hold(negedge G &&& Mux21DTITE_, posedge CD, `LD3SHS_CD_G_REM_posedge_negedge, Notifier);

`else

     if (!D && G && TI) (TE -=> QN) = (`LD3SHS_TE_F_QN_R,`LD3SHS_TE_R_QN_F);
     if (D && G && !TI) (TE +=> QN) = (`LD3SHS_TE_R_QN_R,`LD3SHS_TE_F_QN_F);
      (TI -=> QN) = (`LD3SHS_TI_F_QN_R,`LD3SHS_TI_R_QN_F);
      (D -=> QN) = (`LD3SHS_D_F_QN_R,`LD3SHS_D_R_QN_F);
     if (!D && G && TI) (TE +=> Q) = (`LD3SHS_TE_R_Q_R,`LD3SHS_TE_F_Q_F);
      if (D && G && !TI) (TE -=> Q) = (`LD3SHS_TE_F_Q_R,`LD3SHS_TE_R_Q_F);
      (TI +=> Q) = (`LD3SHS_TI_R_Q_R,`LD3SHS_TI_F_Q_F);
      (D +=> Q) = (`LD3SHS_D_R_Q_R,`LD3SHS_D_F_Q_F);
      (posedge G => (Q +: Mux21DTITE_)) = (`LD3SHS_G_R_Q_R, `LD3SHS_G_R_Q_F);
      (posedge G => (QN -: Mux21DTITE_)) = (`LD3SHS_G_R_QN_R, `LD3SHS_G_R_QN_F);
      (posedge CD => (Q +: 1'b1)) = (`LD3SHS_CD_R_Q_R,`LD3SHS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD3SHS_CD_R_Q_R,`LD3SHS_CD_F_Q_F);
      (posedge CD => (QN +: 1'b0)) = (`LD3SHS_CD_F_QN_R,`LD3SHS_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`LD3SHS_CD_F_QN_R,`LD3SHS_CD_R_QN_F);
 
        $setuphold(negedge G &&& AndXorDTI_CD_, posedge TE, `LD3SHS_TE_G_SETUP_posedge_negedge, `LD3SHS_TE_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& AndXorDTI_CD_, negedge TE, `LD3SHS_TE_G_SETUP_negedge_negedge, `LD3SHS_TE_G_HOLD_negedge_negedge, Notifier);
 
        $setuphold(negedge G &&& AndCDTE_, posedge TI, `LD3SHS_TI_G_SETUP_posedge_negedge, `LD3SHS_TI_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& AndCDTE_, negedge TI, `LD3SHS_TI_G_SETUP_negedge_negedge, `LD3SHS_TI_G_HOLD_negedge_negedge, Notifier);
 
        $setuphold(negedge G &&& AndCDTEX_, posedge D, `LD3SHS_D_G_SETUP_posedge_negedge, `LD3SHS_D_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& AndCDTEX_, negedge D, `LD3SHS_D_G_SETUP_negedge_negedge, `LD3SHS_D_G_HOLD_negedge_negedge, Notifier);
 
      $width(posedge G, `LD3SHS_G_PWH, 0, Notifier);
      $width(negedge CD, `LD3SHS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, negedge G &&& Mux21DTITE_, `LD3SHS_CD_G_REC_posedge_negedge, Notifier);
 
        $hold(negedge G &&& Mux21DTITE_, posedge CD, `LD3SHS_CD_G_REM_posedge_negedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD3SHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:10 and Version :1.1 //
 
//  START 
// CELL LD3SHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD3SHSP_TE_F_QN_R 0.1
`define LD3SHSP_TE_R_QN_F 0.1
`define LD3SHSP_TE_F_QN_F 0.1
`define LD3SHSP_TE_R_QN_R 0.1
`define LD3SHSP_TI_F_QN_R 0.1
`define LD3SHSP_TI_R_QN_F 0.1
`define LD3SHSP_CD_F_QN_R 0.1
`define LD3SHSP_CD_R_QN_F 0.1
`define LD3SHSP_G_R_QN_F 0.1
`define LD3SHSP_G_R_QN_R 0.1
`define LD3SHSP_D_F_QN_R 0.1
`define LD3SHSP_D_R_QN_F 0.1
`define LD3SHSP_TE_F_Q_F 0.1
`define LD3SHSP_TE_R_Q_R 0.1
`define LD3SHSP_TE_F_Q_R 0.1
`define LD3SHSP_TE_R_Q_F 0.1
`define LD3SHSP_TI_F_Q_F 0.1
`define LD3SHSP_TI_R_Q_R 0.1
`define LD3SHSP_CD_F_Q_F 0.1
`define LD3SHSP_CD_R_Q_R 0.1
`define LD3SHSP_G_R_Q_R 0.1
`define LD3SHSP_G_R_Q_F 0.1
`define LD3SHSP_D_F_Q_F 0.1
`define LD3SHSP_D_R_Q_R 0.1
`define LD3SHSP_CD_G_REM_posedge_negedge 0.1
`define LD3SHSP_CD_G_REC_posedge_negedge 0.1
`define LD3SHSP_CD_PWL 0.1
`define LD3SHSP_G_PWH 0.1
`define LD3SHSP_D_G_SETUP_posedge_negedge 0.1
`define LD3SHSP_D_G_SETUP_negedge_negedge 0.1
`define LD3SHSP_D_G_HOLD_posedge_negedge 0.1
`define LD3SHSP_D_G_HOLD_negedge_negedge 0.1
`define LD3SHSP_TI_G_SETUP_posedge_negedge 0.1
`define LD3SHSP_TI_G_SETUP_negedge_negedge 0.1
`define LD3SHSP_TI_G_HOLD_posedge_negedge 0.1
`define LD3SHSP_TI_G_HOLD_negedge_negedge 0.1
`define LD3SHSP_TE_G_SETUP_posedge_negedge 0.1
`define LD3SHSP_TE_G_SETUP_negedge_negedge 0.1
`define LD3SHSP_TE_G_HOLD_posedge_negedge 0.1
`define LD3SHSP_TE_G_HOLD_negedge_negedge 0.1

module LD3SHSP (Q, QN, D, G, CD, TI, TE);

   output Q;
   output QN;
   input D;
   input G;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_LD_P_RN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, G, CD, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   not  (GX, G);
   not  (TEX, TE);
   and  (AndCDTEX_, CD, TEX);
   and  (AndCDTE_, CD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   specify
`ifdef verifault
      if (!D && G && TI) (TE -=> QN) = (`LD3SHSP_TE_F_QN_R,`LD3SHSP_TE_R_QN_F);
      if (D && G && !TI) (TE +=> QN) = (`LD3SHSP_TE_R_QN_R,`LD3SHSP_TE_F_QN_F);
      if (G && CD && TE) (TI -=> QN) = (`LD3SHSP_TI_F_QN_R,`LD3SHSP_TI_R_QN_F);
      if (G && CD && !TE) (D -=> QN) = (`LD3SHSP_D_F_QN_R,`LD3SHSP_D_R_QN_F);
      if (!D && G && TI) (TE +=> Q) = (`LD3SHSP_TE_R_Q_R,`LD3SHSP_TE_F_Q_F);
      if (D && G && !TI) (TE -=> Q) = (`LD3SHSP_TE_F_Q_R,`LD3SHSP_TE_R_Q_F);
      if (G && CD && TE) (TI +=> Q) = (`LD3SHSP_TI_R_Q_R,`LD3SHSP_TI_F_Q_F);
      if (G && CD && !TE) (D +=> Q) = (`LD3SHSP_D_R_Q_R,`LD3SHSP_D_F_Q_F);
      if(!TE) (posedge G => (Q +: D)) = (`LD3SHSP_G_R_Q_R, `LD3SHSP_G_R_Q_F);
      if(TE) (posedge G => (Q +: TI)) = (`LD3SHSP_G_R_Q_R, `LD3SHSP_G_R_Q_F);
      if(!D && TI) (posedge G => (Q +: TE)) = (`LD3SHSP_G_R_Q_R, `LD3SHSP_G_R_Q_F);
      if(!TI && D) (posedge G => (Q -: TE)) = (`LD3SHSP_G_R_Q_R, `LD3SHSP_G_R_Q_F);
      if(!TE) (posedge G => (QN -: D)) = (`LD3SHSP_G_R_QN_R, `LD3SHSP_G_R_QN_F);
      if(TE) (posedge G => (QN -: TI)) = (`LD3SHSP_G_R_QN_R, `LD3SHSP_G_R_QN_F);
      if(!D && TI) (posedge G => (QN -: TE)) = (`LD3SHSP_G_R_QN_R, `LD3SHSP_G_R_QN_F);
      if(!TI && D) (posedge G => (QN +: TE)) = (`LD3SHSP_G_R_QN_R, `LD3SHSP_G_R_QN_F);
      if(D && G && !TE || G && TI && TE) (posedge CD => (Q +: 1'b1)) = (`LD3SHSP_CD_R_Q_R,`LD3SHSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD3SHSP_CD_R_Q_R,`LD3SHSP_CD_F_Q_F);
      if(D && G && !TE || G && TI && TE) (posedge CD => (QN +: 1'b0)) = (`LD3SHSP_CD_F_QN_R,`LD3SHSP_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`LD3SHSP_CD_F_QN_R,`LD3SHSP_CD_R_QN_F);

	$setuphold(negedge G &&& AndXorDTI_CD_, posedge TE, `LD3SHSP_TE_G_SETUP_posedge_negedge, `LD3SHSP_TE_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& AndXorDTI_CD_, negedge TE, `LD3SHSP_TE_G_SETUP_negedge_negedge, `LD3SHSP_TE_G_HOLD_negedge_negedge, Notifier);

	$setuphold(negedge G &&& AndCDTE_, posedge TI, `LD3SHSP_TI_G_SETUP_posedge_negedge, `LD3SHSP_TI_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& AndCDTE_, negedge TI, `LD3SHSP_TI_G_SETUP_negedge_negedge, `LD3SHSP_TI_G_HOLD_negedge_negedge, Notifier);

	$setuphold(negedge G &&& AndCDTEX_, posedge D, `LD3SHSP_D_G_SETUP_posedge_negedge, `LD3SHSP_D_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& AndCDTEX_, negedge D, `LD3SHSP_D_G_SETUP_negedge_negedge, `LD3SHSP_D_G_HOLD_negedge_negedge, Notifier);

      $width(posedge G, `LD3SHSP_G_PWH, 0, Notifier);
      $width(negedge CD, `LD3SHSP_CD_PWL, 0, Notifier);
	$recovery(posedge CD, negedge G &&& Mux21DTITE_, `LD3SHSP_CD_G_REC_posedge_negedge, Notifier);

	$hold(negedge G &&& Mux21DTITE_, posedge CD, `LD3SHSP_CD_G_REM_posedge_negedge, Notifier);

`else

     if (!D && G && TI) (TE -=> QN) = (`LD3SHSP_TE_F_QN_R,`LD3SHSP_TE_R_QN_F);
     if (D && G && !TI) (TE +=> QN) = (`LD3SHSP_TE_R_QN_R,`LD3SHSP_TE_F_QN_F);
      (TI -=> QN) = (`LD3SHSP_TI_F_QN_R,`LD3SHSP_TI_R_QN_F);
      (D -=> QN) = (`LD3SHSP_D_F_QN_R,`LD3SHSP_D_R_QN_F);
     if (!D && G && TI) (TE +=> Q) = (`LD3SHSP_TE_R_Q_R,`LD3SHSP_TE_F_Q_F);
      if (D && G && !TI) (TE -=> Q) = (`LD3SHSP_TE_F_Q_R,`LD3SHSP_TE_R_Q_F);
      (TI +=> Q) = (`LD3SHSP_TI_R_Q_R,`LD3SHSP_TI_F_Q_F);
      (D +=> Q) = (`LD3SHSP_D_R_Q_R,`LD3SHSP_D_F_Q_F);
      (posedge G => (Q +: Mux21DTITE_)) = (`LD3SHSP_G_R_Q_R, `LD3SHSP_G_R_Q_F);
      (posedge G => (QN -: Mux21DTITE_)) = (`LD3SHSP_G_R_QN_R, `LD3SHSP_G_R_QN_F);
      (posedge CD => (Q +: 1'b1)) = (`LD3SHSP_CD_R_Q_R,`LD3SHSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD3SHSP_CD_R_Q_R,`LD3SHSP_CD_F_Q_F);
      (posedge CD => (QN +: 1'b0)) = (`LD3SHSP_CD_F_QN_R,`LD3SHSP_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`LD3SHSP_CD_F_QN_R,`LD3SHSP_CD_R_QN_F);
 
        $setuphold(negedge G &&& AndXorDTI_CD_, posedge TE, `LD3SHSP_TE_G_SETUP_posedge_negedge, `LD3SHSP_TE_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& AndXorDTI_CD_, negedge TE, `LD3SHSP_TE_G_SETUP_negedge_negedge, `LD3SHSP_TE_G_HOLD_negedge_negedge, Notifier);
 
        $setuphold(negedge G &&& AndCDTE_, posedge TI, `LD3SHSP_TI_G_SETUP_posedge_negedge, `LD3SHSP_TI_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& AndCDTE_, negedge TI, `LD3SHSP_TI_G_SETUP_negedge_negedge, `LD3SHSP_TI_G_HOLD_negedge_negedge, Notifier);
 
        $setuphold(negedge G &&& AndCDTEX_, posedge D, `LD3SHSP_D_G_SETUP_posedge_negedge, `LD3SHSP_D_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& AndCDTEX_, negedge D, `LD3SHSP_D_G_SETUP_negedge_negedge, `LD3SHSP_D_G_HOLD_negedge_negedge, Notifier);
 
      $width(posedge G, `LD3SHSP_G_PWH, 0, Notifier);
      $width(negedge CD, `LD3SHSP_CD_PWL, 0, Notifier);
        $recovery(posedge CD, negedge G &&& Mux21DTITE_, `LD3SHSP_CD_G_REC_posedge_negedge, Notifier);
 
        $hold(negedge G &&& Mux21DTITE_, posedge CD, `LD3SHSP_CD_G_REM_posedge_negedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD3SHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:10 and Version :1.1 //
 
//  START 
// CELL LD3SQHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD3SQHS_TE_F_Q_F 0.1
`define LD3SQHS_TE_R_Q_R 0.1
`define LD3SQHS_TE_F_Q_R 0.1
`define LD3SQHS_TE_R_Q_F 0.1
`define LD3SQHS_TI_F_Q_F 0.1
`define LD3SQHS_TI_R_Q_R 0.1
`define LD3SQHS_CD_F_Q_F 0.1
`define LD3SQHS_CD_R_Q_R 0.1
`define LD3SQHS_G_R_Q_R 0.1
`define LD3SQHS_G_R_Q_F 0.1
`define LD3SQHS_D_F_Q_F 0.1
`define LD3SQHS_D_R_Q_R 0.1
`define LD3SQHS_TE_G_HOLD_posedge_negedge 0.1
`define LD3SQHS_TE_G_HOLD_negedge_negedge 0.1
`define LD3SQHS_TE_G_SETUP_posedge_negedge 0.1
`define LD3SQHS_TE_G_SETUP_negedge_negedge 0.1
`define LD3SQHS_TI_G_HOLD_posedge_negedge 0.1
`define LD3SQHS_TI_G_HOLD_negedge_negedge 0.1
`define LD3SQHS_TI_G_SETUP_posedge_negedge 0.1
`define LD3SQHS_TI_G_SETUP_negedge_negedge 0.1
`define LD3SQHS_D_G_HOLD_posedge_negedge 0.1
`define LD3SQHS_D_G_HOLD_negedge_negedge 0.1
`define LD3SQHS_D_G_SETUP_posedge_negedge 0.1
`define LD3SQHS_D_G_SETUP_negedge_negedge 0.1
`define LD3SQHS_G_PWH 0.1
`define LD3SQHS_CD_PWL 0.1
`define LD3SQHS_CD_G_REC_posedge_negedge 0.1
`define LD3SQHS_CD_G_REM_posedge_negedge 0.1

module LD3SQHS (Q, D, G, CD, TI, TE);

   output Q;
   input D;
   input G;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_LD_P_RN_NOTI u1 (IQ, Mux21DTITE_, G, CD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   not  (GX, G);
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);

   specify
`ifdef verifault
      if (!D && G && TI) (TE +=> Q) = (`LD3SQHS_TE_R_Q_R,`LD3SQHS_TE_F_Q_F);
      if (D && G && !TI) (TE -=> Q) = (`LD3SQHS_TE_F_Q_R,`LD3SQHS_TE_R_Q_F);
      if (G && CD && TE) (TI +=> Q) = (`LD3SQHS_TI_R_Q_R,`LD3SQHS_TI_F_Q_F);
      if (G && CD && !TE) (D +=> Q) = (`LD3SQHS_D_R_Q_R,`LD3SQHS_D_F_Q_F);
      if(!TE && CD) (posedge G => (Q +: D)) = (`LD3SQHS_G_R_Q_R, `LD3SQHS_G_R_Q_F);
      if(TE && CD) (posedge G => (Q +: TI)) = (`LD3SQHS_G_R_Q_R, `LD3SQHS_G_R_Q_F);
      if(!D && TI && CD) (posedge G => (Q +: TE)) = (`LD3SQHS_G_R_Q_R, `LD3SQHS_G_R_Q_F);
      if(!TI && D && CD) (posedge G => (Q -: TE)) = (`LD3SQHS_G_R_Q_R, `LD3SQHS_G_R_Q_F);
      if(D && G && !TE || G && TI && TE) (posedge CD => (Q +: 1'b1)) = (`LD3SQHS_CD_R_Q_R,`LD3SQHS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD3SQHS_CD_R_Q_R,`LD3SQHS_CD_F_Q_F);

	$setuphold(negedge G &&& AndXorDTI_CD_, posedge TE, `LD3SQHS_TE_G_SETUP_posedge_negedge, `LD3SQHS_TE_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& AndXorDTI_CD_, negedge TE, `LD3SQHS_TE_G_SETUP_negedge_negedge, `LD3SQHS_TE_G_HOLD_negedge_negedge, Notifier);

	$setuphold(negedge G &&& AndCDTE_, posedge TI, `LD3SQHS_TI_G_SETUP_posedge_negedge, `LD3SQHS_TI_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& AndCDTE_, negedge TI, `LD3SQHS_TI_G_SETUP_negedge_negedge, `LD3SQHS_TI_G_HOLD_negedge_negedge, Notifier);

	$setuphold(negedge G &&& AndCDTEX_, posedge D, `LD3SQHS_D_G_SETUP_posedge_negedge, `LD3SQHS_D_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& AndCDTEX_, negedge D, `LD3SQHS_D_G_SETUP_negedge_negedge, `LD3SQHS_D_G_HOLD_negedge_negedge, Notifier);

      $width(posedge G, `LD3SQHS_G_PWH, 0, Notifier);
      $width(negedge CD, `LD3SQHS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, negedge G &&& Mux21DTITE_, `LD3SQHS_CD_G_REC_posedge_negedge, Notifier);

	$hold(negedge G &&& Mux21DTITE_, posedge CD, `LD3SQHS_CD_G_REM_posedge_negedge, Notifier);

`else
      if (!D && G && TI) (TE +=> Q) = (`LD3SQHS_TE_R_Q_R,`LD3SQHS_TE_F_Q_F);
      if (D && G && !TI) (TE -=> Q) = (`LD3SQHS_TE_F_Q_R,`LD3SQHS_TE_R_Q_F);
      (TI +=> Q) = (`LD3SQHS_TI_R_Q_R,`LD3SQHS_TI_F_Q_F);
      (D +=> Q) = (`LD3SQHS_D_R_Q_R,`LD3SQHS_D_F_Q_F);
      (posedge G => (Q +: Mux21DTITE_)) = (`LD3SQHS_G_R_Q_R, `LD3SQHS_G_R_Q_F);
      (posedge CD => (Q +: 1'b1)) = (`LD3SQHS_CD_R_Q_R,`LD3SQHS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD3SQHS_CD_R_Q_R,`LD3SQHS_CD_F_Q_F);
 
        $setuphold(negedge G &&& AndXorDTI_CD_, posedge TE, `LD3SQHS_TE_G_SETUP_posedge_negedge, `LD3SQHS_TE_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& AndXorDTI_CD_, negedge TE, `LD3SQHS_TE_G_SETUP_negedge_negedge, `LD3SQHS_TE_G_HOLD_negedge_negedge, Notifier);
 
        $setuphold(negedge G &&& AndCDTE_, posedge TI, `LD3SQHS_TI_G_SETUP_posedge_negedge, `LD3SQHS_TI_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& AndCDTE_, negedge TI, `LD3SQHS_TI_G_SETUP_negedge_negedge, `LD3SQHS_TI_G_HOLD_negedge_negedge, Notifier);
 
        $setuphold(negedge G &&& AndCDTEX_, posedge D, `LD3SQHS_D_G_SETUP_posedge_negedge, `LD3SQHS_D_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& AndCDTEX_, negedge D, `LD3SQHS_D_G_SETUP_negedge_negedge, `LD3SQHS_D_G_HOLD_negedge_negedge, Notifier);
 
      $width(posedge G, `LD3SQHS_G_PWH, 0, Notifier);
      $width(negedge CD, `LD3SQHS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, negedge G &&& Mux21DTITE_, `LD3SQHS_CD_G_REC_posedge_negedge, Notifier);
 
        $hold(negedge G &&& Mux21DTITE_, posedge CD, `LD3SQHS_CD_G_REM_posedge_negedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD3SQHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:10 and Version :1.1 //
 
//  START 
// CELL LD3SQHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD3SQHSP_TE_F_Q_F 0.1
`define LD3SQHSP_TE_R_Q_R 0.1
`define LD3SQHSP_TE_F_Q_R 0.1
`define LD3SQHSP_TE_R_Q_F 0.1
`define LD3SQHSP_TI_F_Q_F 0.1
`define LD3SQHSP_TI_R_Q_R 0.1
`define LD3SQHSP_CD_F_Q_F 0.1
`define LD3SQHSP_CD_R_Q_R 0.1
`define LD3SQHSP_G_R_Q_R 0.1
`define LD3SQHSP_G_R_Q_F 0.1
`define LD3SQHSP_D_F_Q_F 0.1
`define LD3SQHSP_D_R_Q_R 0.1
`define LD3SQHSP_TE_G_HOLD_posedge_negedge 0.1
`define LD3SQHSP_TE_G_HOLD_negedge_negedge 0.1
`define LD3SQHSP_TE_G_SETUP_posedge_negedge 0.1
`define LD3SQHSP_TE_G_SETUP_negedge_negedge 0.1
`define LD3SQHSP_TI_G_HOLD_posedge_negedge 0.1
`define LD3SQHSP_TI_G_HOLD_negedge_negedge 0.1
`define LD3SQHSP_TI_G_SETUP_posedge_negedge 0.1
`define LD3SQHSP_TI_G_SETUP_negedge_negedge 0.1
`define LD3SQHSP_D_G_HOLD_posedge_negedge 0.1
`define LD3SQHSP_D_G_HOLD_negedge_negedge 0.1
`define LD3SQHSP_D_G_SETUP_posedge_negedge 0.1
`define LD3SQHSP_D_G_SETUP_negedge_negedge 0.1
`define LD3SQHSP_G_PWH 0.1
`define LD3SQHSP_CD_PWL 0.1
`define LD3SQHSP_CD_G_REC_posedge_negedge 0.1
`define LD3SQHSP_CD_G_REM_posedge_negedge 0.1

module LD3SQHSP (Q, D, G, CD, TI, TE);

   output Q;
   input D;
   input G;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_LD_P_RN_NOTI u1 (IQ, Mux21DTITE_, G, CD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   not  (GX, G);
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);

   specify
`ifdef verifault
      if (!D && G && TI) (TE +=> Q) = (`LD3SQHSP_TE_R_Q_R,`LD3SQHSP_TE_F_Q_F);
      if (D && G && !TI) (TE -=> Q) = (`LD3SQHSP_TE_F_Q_R,`LD3SQHSP_TE_R_Q_F);
      if (G && CD && TE) (TI +=> Q) = (`LD3SQHSP_TI_R_Q_R,`LD3SQHSP_TI_F_Q_F);
      if (G && CD && !TE) (D +=> Q) = (`LD3SQHSP_D_R_Q_R,`LD3SQHSP_D_F_Q_F);
      if(!TE && CD) (posedge G => (Q +: D)) = (`LD3SQHSP_G_R_Q_R, `LD3SQHSP_G_R_Q_F);
      if(TE && CD) (posedge G => (Q +: TI)) = (`LD3SQHSP_G_R_Q_R, `LD3SQHSP_G_R_Q_F);
      if(!D && TI && CD) (posedge G => (Q +: TE)) = (`LD3SQHSP_G_R_Q_R, `LD3SQHSP_G_R_Q_F);
      if(!TI && D && CD) (posedge G => (Q -: TE)) = (`LD3SQHSP_G_R_Q_R, `LD3SQHSP_G_R_Q_F);
      if(D && G && !TE || G && TI && TE) (posedge CD => (Q +: 1'b1)) = (`LD3SQHSP_CD_R_Q_R,`LD3SQHSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD3SQHSP_CD_R_Q_R,`LD3SQHSP_CD_F_Q_F);

	$setuphold(negedge G &&& AndXorDTI_CD_, posedge TE, `LD3SQHSP_TE_G_SETUP_posedge_negedge, `LD3SQHSP_TE_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& AndXorDTI_CD_, negedge TE, `LD3SQHSP_TE_G_SETUP_negedge_negedge, `LD3SQHSP_TE_G_HOLD_negedge_negedge, Notifier);

	$setuphold(negedge G &&& AndCDTE_, posedge TI, `LD3SQHSP_TI_G_SETUP_posedge_negedge, `LD3SQHSP_TI_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& AndCDTE_, negedge TI, `LD3SQHSP_TI_G_SETUP_negedge_negedge, `LD3SQHSP_TI_G_HOLD_negedge_negedge, Notifier);

	$setuphold(negedge G &&& AndCDTEX_, posedge D, `LD3SQHSP_D_G_SETUP_posedge_negedge, `LD3SQHSP_D_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& AndCDTEX_, negedge D, `LD3SQHSP_D_G_SETUP_negedge_negedge, `LD3SQHSP_D_G_HOLD_negedge_negedge, Notifier);

      $width(posedge G, `LD3SQHSP_G_PWH, 0, Notifier);
      $width(negedge CD, `LD3SQHSP_CD_PWL, 0, Notifier);
	$recovery(posedge CD, negedge G &&& Mux21DTITE_, `LD3SQHSP_CD_G_REC_posedge_negedge, Notifier);

	$hold(negedge G &&& Mux21DTITE_, posedge CD, `LD3SQHSP_CD_G_REM_posedge_negedge, Notifier);

`else
      if (!D && G && TI) (TE +=> Q) = (`LD3SQHSP_TE_R_Q_R,`LD3SQHSP_TE_F_Q_F);
      if (D && G && !TI) (TE -=> Q) = (`LD3SQHSP_TE_F_Q_R,`LD3SQHSP_TE_R_Q_F);
      (TI +=> Q) = (`LD3SQHSP_TI_R_Q_R,`LD3SQHSP_TI_F_Q_F);
      (D +=> Q) = (`LD3SQHSP_D_R_Q_R,`LD3SQHSP_D_F_Q_F);
      (posedge G => (Q +: Mux21DTITE_)) = (`LD3SQHSP_G_R_Q_R, `LD3SQHSP_G_R_Q_F);
      (posedge CD => (Q +: 1'b1)) = (`LD3SQHSP_CD_R_Q_R,`LD3SQHSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD3SQHSP_CD_R_Q_R,`LD3SQHSP_CD_F_Q_F);
 
        $setuphold(negedge G &&& AndXorDTI_CD_, posedge TE, `LD3SQHSP_TE_G_SETUP_posedge_negedge, `LD3SQHSP_TE_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& AndXorDTI_CD_, negedge TE, `LD3SQHSP_TE_G_SETUP_negedge_negedge, `LD3SQHSP_TE_G_HOLD_negedge_negedge, Notifier);
 
        $setuphold(negedge G &&& AndCDTE_, posedge TI, `LD3SQHSP_TI_G_SETUP_posedge_negedge, `LD3SQHSP_TI_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& AndCDTE_, negedge TI, `LD3SQHSP_TI_G_SETUP_negedge_negedge, `LD3SQHSP_TI_G_HOLD_negedge_negedge, Notifier);
 
        $setuphold(negedge G &&& AndCDTEX_, posedge D, `LD3SQHSP_D_G_SETUP_posedge_negedge, `LD3SQHSP_D_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& AndCDTEX_, negedge D, `LD3SQHSP_D_G_SETUP_negedge_negedge, `LD3SQHSP_D_G_HOLD_negedge_negedge, Notifier);
 
      $width(posedge G, `LD3SQHSP_G_PWH, 0, Notifier);
      $width(negedge CD, `LD3SQHSP_CD_PWL, 0, Notifier);
        $recovery(posedge CD, negedge G &&& Mux21DTITE_, `LD3SQHSP_CD_G_REC_posedge_negedge, Notifier);
 
        $hold(negedge G &&& Mux21DTITE_, posedge CD, `LD3SQHSP_CD_G_REM_posedge_negedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD3SQHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:10 and Version :1.1 //
 
//  START 
// CELL LD3SQHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD3SQHSX4_TE_F_Q_F 0.1
`define LD3SQHSX4_TE_R_Q_R 0.1
`define LD3SQHSX4_TE_F_Q_R 0.1
`define LD3SQHSX4_TE_R_Q_F 0.1
`define LD3SQHSX4_TI_F_Q_F 0.1
`define LD3SQHSX4_TI_R_Q_R 0.1
`define LD3SQHSX4_CD_F_Q_F 0.1
`define LD3SQHSX4_CD_R_Q_R 0.1
`define LD3SQHSX4_G_R_Q_R 0.1
`define LD3SQHSX4_G_R_Q_F 0.1
`define LD3SQHSX4_D_F_Q_F 0.1
`define LD3SQHSX4_D_R_Q_R 0.1
`define LD3SQHSX4_TE_G_HOLD_posedge_negedge 0.1
`define LD3SQHSX4_TE_G_HOLD_negedge_negedge 0.1
`define LD3SQHSX4_TE_G_SETUP_posedge_negedge 0.1
`define LD3SQHSX4_TE_G_SETUP_negedge_negedge 0.1
`define LD3SQHSX4_TI_G_HOLD_posedge_negedge 0.1
`define LD3SQHSX4_TI_G_HOLD_negedge_negedge 0.1
`define LD3SQHSX4_TI_G_SETUP_posedge_negedge 0.1
`define LD3SQHSX4_TI_G_SETUP_negedge_negedge 0.1
`define LD3SQHSX4_D_G_HOLD_posedge_negedge 0.1
`define LD3SQHSX4_D_G_HOLD_negedge_negedge 0.1
`define LD3SQHSX4_D_G_SETUP_posedge_negedge 0.1
`define LD3SQHSX4_D_G_SETUP_negedge_negedge 0.1
`define LD3SQHSX4_G_PWH 0.1
`define LD3SQHSX4_CD_PWL 0.1
`define LD3SQHSX4_CD_G_REC_posedge_negedge 0.1
`define LD3SQHSX4_CD_G_REM_posedge_negedge 0.1

module LD3SQHSX4 (Q, D, G, CD, TI, TE);

   output Q;
   input D;
   input G;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_LD_P_RN_NOTI u1 (IQ, Mux21DTITE_, G, CD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   not  (GX, G);
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);

   specify
`ifdef verifault
      if (!D && G && TI) (TE +=> Q) = (`LD3SQHSX4_TE_R_Q_R,`LD3SQHSX4_TE_F_Q_F);
      if (D && G && !TI) (TE -=> Q) = (`LD3SQHSX4_TE_F_Q_R,`LD3SQHSX4_TE_R_Q_F);
      if (G && CD && TE) (TI +=> Q) = (`LD3SQHSX4_TI_R_Q_R,`LD3SQHSX4_TI_F_Q_F);
      if (G && CD && !TE) (D +=> Q) = (`LD3SQHSX4_D_R_Q_R,`LD3SQHSX4_D_F_Q_F);
      if(!TE && CD) (posedge G => (Q +: D)) = (`LD3SQHSX4_G_R_Q_R, `LD3SQHSX4_G_R_Q_F);
      if(TE && CD) (posedge G => (Q +: TI)) = (`LD3SQHSX4_G_R_Q_R, `LD3SQHSX4_G_R_Q_F);
      if(!D && TI && CD) (posedge G => (Q +: TE)) = (`LD3SQHSX4_G_R_Q_R, `LD3SQHSX4_G_R_Q_F);
      if(!TI && D && CD) (posedge G => (Q -: TE)) = (`LD3SQHSX4_G_R_Q_R, `LD3SQHSX4_G_R_Q_F);
      if(D && G && !TE || G && TI && TE) (posedge CD => (Q +: 1'b1)) = (`LD3SQHSX4_CD_R_Q_R,`LD3SQHSX4_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD3SQHSX4_CD_R_Q_R,`LD3SQHSX4_CD_F_Q_F);

	$setuphold(negedge G &&& AndXorDTI_CD_, posedge TE, `LD3SQHSX4_TE_G_SETUP_posedge_negedge, `LD3SQHSX4_TE_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& AndXorDTI_CD_, negedge TE, `LD3SQHSX4_TE_G_SETUP_negedge_negedge, `LD3SQHSX4_TE_G_HOLD_negedge_negedge, Notifier);

	$setuphold(negedge G &&& AndCDTE_, posedge TI, `LD3SQHSX4_TI_G_SETUP_posedge_negedge, `LD3SQHSX4_TI_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& AndCDTE_, negedge TI, `LD3SQHSX4_TI_G_SETUP_negedge_negedge, `LD3SQHSX4_TI_G_HOLD_negedge_negedge, Notifier);

	$setuphold(negedge G &&& AndCDTEX_, posedge D, `LD3SQHSX4_D_G_SETUP_posedge_negedge, `LD3SQHSX4_D_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& AndCDTEX_, negedge D, `LD3SQHSX4_D_G_SETUP_negedge_negedge, `LD3SQHSX4_D_G_HOLD_negedge_negedge, Notifier);

      $width(posedge G, `LD3SQHSX4_G_PWH, 0, Notifier);
      $width(negedge CD, `LD3SQHSX4_CD_PWL, 0, Notifier);
	$recovery(posedge CD, negedge G &&& Mux21DTITE_, `LD3SQHSX4_CD_G_REC_posedge_negedge, Notifier);

	$hold(negedge G &&& Mux21DTITE_, posedge CD, `LD3SQHSX4_CD_G_REM_posedge_negedge, Notifier);

`else
      if (!D && G && TI) (TE +=> Q) = (`LD3SQHSX4_TE_R_Q_R,`LD3SQHSX4_TE_F_Q_F);
      if (D && G && !TI) (TE -=> Q) = (`LD3SQHSX4_TE_F_Q_R,`LD3SQHSX4_TE_R_Q_F);
      (TI +=> Q) = (`LD3SQHSX4_TI_R_Q_R,`LD3SQHSX4_TI_F_Q_F);
      (D +=> Q) = (`LD3SQHSX4_D_R_Q_R,`LD3SQHSX4_D_F_Q_F);
      (posedge G => (Q +: Mux21DTITE_)) = (`LD3SQHSX4_G_R_Q_R, `LD3SQHSX4_G_R_Q_F);
      (posedge CD => (Q +: 1'b1)) = (`LD3SQHSX4_CD_R_Q_R,`LD3SQHSX4_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD3SQHSX4_CD_R_Q_R,`LD3SQHSX4_CD_F_Q_F);
 
        $setuphold(negedge G &&& AndXorDTI_CD_, posedge TE, `LD3SQHSX4_TE_G_SETUP_posedge_negedge, `LD3SQHSX4_TE_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& AndXorDTI_CD_, negedge TE, `LD3SQHSX4_TE_G_SETUP_negedge_negedge, `LD3SQHSX4_TE_G_HOLD_negedge_negedge, Notifier);
 
        $setuphold(negedge G &&& AndCDTE_, posedge TI, `LD3SQHSX4_TI_G_SETUP_posedge_negedge, `LD3SQHSX4_TI_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& AndCDTE_, negedge TI, `LD3SQHSX4_TI_G_SETUP_negedge_negedge, `LD3SQHSX4_TI_G_HOLD_negedge_negedge, Notifier);
 
        $setuphold(negedge G &&& AndCDTEX_, posedge D, `LD3SQHSX4_D_G_SETUP_posedge_negedge, `LD3SQHSX4_D_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& AndCDTEX_, negedge D, `LD3SQHSX4_D_G_SETUP_negedge_negedge, `LD3SQHSX4_D_G_HOLD_negedge_negedge, Notifier);
 
      $width(posedge G, `LD3SQHSX4_G_PWH, 0, Notifier);
      $width(negedge CD, `LD3SQHSX4_CD_PWL, 0, Notifier);
        $recovery(posedge CD, negedge G &&& Mux21DTITE_, `LD3SQHSX4_CD_G_REC_posedge_negedge, Notifier);
 
        $hold(negedge G &&& Mux21DTITE_, posedge CD, `LD3SQHSX4_CD_G_REM_posedge_negedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD3SQHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:10 and Version :1.1 //
 
//  START 
// CELL LD4HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD4HS_CD_F_QN_R 0.1
`define LD4HS_CD_R_QN_F 0.1
`define LD4HS_GN_F_QN_F 0.1
`define LD4HS_GN_F_QN_R 0.1
`define LD4HS_D_F_QN_R 0.1
`define LD4HS_D_R_QN_F 0.1
`define LD4HS_CD_F_Q_F 0.1
`define LD4HS_CD_R_Q_R 0.1
`define LD4HS_GN_F_Q_R 0.1
`define LD4HS_GN_F_Q_F 0.1
`define LD4HS_D_F_Q_F 0.1
`define LD4HS_D_R_Q_R 0.1
`define LD4HS_CD_GN_REM_posedge_posedge 0.1
`define LD4HS_CD_GN_REC_posedge_posedge 0.1
`define LD4HS_CD_PWL 0.1
`define LD4HS_GN_PWL 0.1
`define LD4HS_D_GN_SETUP_posedge_posedge 0.1
`define LD4HS_D_GN_SETUP_negedge_posedge 0.1
`define LD4HS_D_GN_HOLD_posedge_posedge 0.1
`define LD4HS_D_GN_HOLD_negedge_posedge 0.1

module LD4HS (Q, QN, D, GN, CD);

   output Q;
   output QN;
   input D;
   input GN;
   input CD;


   reg Notifier;


   U_LD_N_RN_NOTI u0 (   // Verilog Seq UDP
      IQ, D, GN, CD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if (!GN && CD) (D -=> QN) = (`LD4HS_D_F_QN_R,`LD4HS_D_R_QN_F);
      if (!GN && CD) (D +=> Q) = (`LD4HS_D_R_Q_R,`LD4HS_D_F_Q_F);
      (negedge GN => (Q +: D)) = (`LD4HS_GN_F_Q_R, `LD4HS_GN_F_Q_F);
      (negedge GN => (QN -: D)) = (`LD4HS_GN_F_QN_R, `LD4HS_GN_F_QN_F);
      if(D && !GN) (posedge CD => (Q +: 1'b1)) = (`LD4HS_CD_R_Q_R,`LD4HS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD4HS_CD_R_Q_R,`LD4HS_CD_F_Q_F);
      if(D && !GN) (posedge CD => (QN +: 1'b0)) = (`LD4HS_CD_F_QN_R,`LD4HS_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`LD4HS_CD_F_QN_R,`LD4HS_CD_R_QN_F);

	$setuphold(posedge GN &&& CD, posedge D, `LD4HS_D_GN_SETUP_posedge_posedge, `LD4HS_D_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& CD, negedge D, `LD4HS_D_GN_SETUP_negedge_posedge, `LD4HS_D_GN_HOLD_negedge_posedge, Notifier);

      $width(negedge GN, `LD4HS_GN_PWL, 0, Notifier);
      $width(negedge CD, `LD4HS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge GN &&& D, `LD4HS_CD_GN_REC_posedge_posedge, Notifier);

	$hold(posedge GN &&& D, posedge CD, `LD4HS_CD_GN_REM_posedge_posedge, Notifier);

`else


      (D -=> QN) = (`LD4HS_D_F_QN_R,`LD4HS_D_R_QN_F);
      (D +=> Q) = (`LD4HS_D_R_Q_R,`LD4HS_D_F_Q_F);
      (negedge GN => (Q +: D)) = (`LD4HS_GN_F_Q_R, `LD4HS_GN_F_Q_F);
      (negedge GN => (QN -: D)) = (`LD4HS_GN_F_QN_R, `LD4HS_GN_F_QN_F);
      (posedge CD => (Q +: 1'b1)) = (`LD4HS_CD_R_Q_R,`LD4HS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD4HS_CD_R_Q_R,`LD4HS_CD_F_Q_F);
      (posedge CD => (QN +: 1'b0)) = (`LD4HS_CD_F_QN_R,`LD4HS_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`LD4HS_CD_F_QN_R,`LD4HS_CD_R_QN_F);
 
        $setuphold(posedge GN &&& CD, posedge D, `LD4HS_D_GN_SETUP_posedge_posedge, `LD4HS_D_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& CD, negedge D, `LD4HS_D_GN_SETUP_negedge_posedge, `LD4HS_D_GN_HOLD_negedge_posedge, Notifier);
 
      $width(negedge GN, `LD4HS_GN_PWL, 0, Notifier);
      $width(negedge CD, `LD4HS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge GN &&& D, `LD4HS_CD_GN_REC_posedge_posedge, Notifier);
 
        $hold(posedge GN &&& D, posedge CD, `LD4HS_CD_GN_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD4HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:17 and Version :1.1 //
 
//  START 
// CELL LD4HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD4HSP_CD_F_QN_R 0.1
`define LD4HSP_CD_R_QN_F 0.1
`define LD4HSP_GN_F_QN_F 0.1
`define LD4HSP_GN_F_QN_R 0.1
`define LD4HSP_D_F_QN_R 0.1
`define LD4HSP_D_R_QN_F 0.1
`define LD4HSP_CD_F_Q_F 0.1
`define LD4HSP_CD_R_Q_R 0.1
`define LD4HSP_GN_F_Q_R 0.1
`define LD4HSP_GN_F_Q_F 0.1
`define LD4HSP_D_F_Q_F 0.1
`define LD4HSP_D_R_Q_R 0.1
`define LD4HSP_CD_GN_REM_posedge_posedge 0.1
`define LD4HSP_CD_GN_REC_posedge_posedge 0.1
`define LD4HSP_CD_PWL 0.1
`define LD4HSP_GN_PWL 0.1
`define LD4HSP_D_GN_SETUP_posedge_posedge 0.1
`define LD4HSP_D_GN_SETUP_negedge_posedge 0.1
`define LD4HSP_D_GN_HOLD_posedge_posedge 0.1
`define LD4HSP_D_GN_HOLD_negedge_posedge 0.1

module LD4HSP (Q, QN, D, GN, CD);

   output Q;
   output QN;
   input D;
   input GN;
   input CD;


   reg Notifier;


   U_LD_N_RN_NOTI u0 (   // Verilog Seq UDP
      IQ, D, GN, CD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if (!GN && CD) (D -=> QN) = (`LD4HSP_D_F_QN_R,`LD4HSP_D_R_QN_F);
      if (!GN && CD) (D +=> Q) = (`LD4HSP_D_R_Q_R,`LD4HSP_D_F_Q_F);
      (negedge GN => (Q +: D)) = (`LD4HSP_GN_F_Q_R, `LD4HSP_GN_F_Q_F);
      (negedge GN => (QN -: D)) = (`LD4HSP_GN_F_QN_R, `LD4HSP_GN_F_QN_F);
      if(D && !GN) (posedge CD => (Q +: 1'b1)) = (`LD4HSP_CD_R_Q_R,`LD4HSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD4HSP_CD_R_Q_R,`LD4HSP_CD_F_Q_F);
      if(D && !GN) (posedge CD => (QN +: 1'b0)) = (`LD4HSP_CD_F_QN_R,`LD4HSP_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`LD4HSP_CD_F_QN_R,`LD4HSP_CD_R_QN_F);

	$setuphold(posedge GN &&& CD, posedge D, `LD4HSP_D_GN_SETUP_posedge_posedge, `LD4HSP_D_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& CD, negedge D, `LD4HSP_D_GN_SETUP_negedge_posedge, `LD4HSP_D_GN_HOLD_negedge_posedge, Notifier);

      $width(negedge GN, `LD4HSP_GN_PWL, 0, Notifier);
      $width(negedge CD, `LD4HSP_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge GN &&& D, `LD4HSP_CD_GN_REC_posedge_posedge, Notifier);

	$hold(posedge GN &&& D, posedge CD, `LD4HSP_CD_GN_REM_posedge_posedge, Notifier);

`else


      (D -=> QN) = (`LD4HSP_D_F_QN_R,`LD4HSP_D_R_QN_F);
      (D +=> Q) = (`LD4HSP_D_R_Q_R,`LD4HSP_D_F_Q_F);
      (negedge GN => (Q +: D)) = (`LD4HSP_GN_F_Q_R, `LD4HSP_GN_F_Q_F);
      (negedge GN => (QN -: D)) = (`LD4HSP_GN_F_QN_R, `LD4HSP_GN_F_QN_F);
      (posedge CD => (Q +: 1'b1)) = (`LD4HSP_CD_R_Q_R,`LD4HSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD4HSP_CD_R_Q_R,`LD4HSP_CD_F_Q_F);
      (posedge CD => (QN +: 1'b0)) = (`LD4HSP_CD_F_QN_R,`LD4HSP_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`LD4HSP_CD_F_QN_R,`LD4HSP_CD_R_QN_F);
 
        $setuphold(posedge GN &&& CD, posedge D, `LD4HSP_D_GN_SETUP_posedge_posedge, `LD4HSP_D_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& CD, negedge D, `LD4HSP_D_GN_SETUP_negedge_posedge, `LD4HSP_D_GN_HOLD_negedge_posedge, Notifier);
 
      $width(negedge GN, `LD4HSP_GN_PWL, 0, Notifier);
      $width(negedge CD, `LD4HSP_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge GN &&& D, `LD4HSP_CD_GN_REC_posedge_posedge, Notifier);
 
        $hold(posedge GN &&& D, posedge CD, `LD4HSP_CD_GN_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD4HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:17 and Version :1.1 //
 
//  START 
// CELL LD4QHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD4QHS_CD_F_Q_F 0.1
`define LD4QHS_CD_R_Q_R 0.1
`define LD4QHS_GN_F_Q_R 0.1
`define LD4QHS_GN_F_Q_F 0.1
`define LD4QHS_D_F_Q_F 0.1
`define LD4QHS_D_R_Q_R 0.1
`define LD4QHS_D_GN_HOLD_posedge_posedge 0.1
`define LD4QHS_D_GN_HOLD_negedge_posedge 0.1
`define LD4QHS_D_GN_SETUP_posedge_posedge 0.1
`define LD4QHS_D_GN_SETUP_negedge_posedge 0.1
`define LD4QHS_GN_PWL 0.1
`define LD4QHS_CD_PWL 0.1
`define LD4QHS_CD_GN_REC_posedge_posedge 0.1
`define LD4QHS_CD_GN_REM_posedge_posedge 0.1

module LD4QHS (Q, D, GN, CD);

   output Q;
   input D;
   input GN;
   input CD;


   reg Notifier;


   U_LD_N_RN_NOTI u0 (IQ, D, GN, CD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if (!GN && CD) (D +=> Q) = (`LD4QHS_D_R_Q_R,`LD4QHS_D_F_Q_F);
      if(CD) (negedge GN => (Q +: D)) = (`LD4QHS_GN_F_Q_R, `LD4QHS_GN_F_Q_F);
      if(D && !GN) (posedge CD => (Q +: 1'b1)) = (`LD4QHS_CD_R_Q_R,`LD4QHS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD4QHS_CD_R_Q_R,`LD4QHS_CD_F_Q_F);

	$setuphold(posedge GN &&& CD, posedge D, `LD4QHS_D_GN_SETUP_posedge_posedge, `LD4QHS_D_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& CD, negedge D, `LD4QHS_D_GN_SETUP_negedge_posedge, `LD4QHS_D_GN_HOLD_negedge_posedge, Notifier);

      $width(negedge GN, `LD4QHS_GN_PWL, 0, Notifier);
      $width(negedge CD, `LD4QHS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge GN &&& D, `LD4QHS_CD_GN_REC_posedge_posedge, Notifier);

	$hold(posedge GN &&& D, posedge CD, `LD4QHS_CD_GN_REM_posedge_posedge, Notifier);

`else

      (D +=> Q) = (`LD4QHS_D_R_Q_R,`LD4QHS_D_F_Q_F);
      (negedge GN => (Q +: D)) = (`LD4QHS_GN_F_Q_R, `LD4QHS_GN_F_Q_F);
      (posedge CD => (Q +: 1'b1)) = (`LD4QHS_CD_R_Q_R,`LD4QHS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD4QHS_CD_R_Q_R,`LD4QHS_CD_F_Q_F);
 
        $setuphold(posedge GN &&& CD, posedge D, `LD4QHS_D_GN_SETUP_posedge_posedge, `LD4QHS_D_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& CD, negedge D, `LD4QHS_D_GN_SETUP_negedge_posedge, `LD4QHS_D_GN_HOLD_negedge_posedge, Notifier);
 
      $width(negedge GN, `LD4QHS_GN_PWL, 0, Notifier);
      $width(negedge CD, `LD4QHS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge GN &&& D, `LD4QHS_CD_GN_REC_posedge_posedge, Notifier);
 
        $hold(posedge GN &&& D, posedge CD, `LD4QHS_CD_GN_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD4QHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:17 and Version :1.1 //
 
//  START 
// CELL LD4QHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD4QHSP_CD_F_Q_F 0.1
`define LD4QHSP_CD_R_Q_R 0.1
`define LD4QHSP_GN_F_Q_R 0.1
`define LD4QHSP_GN_F_Q_F 0.1
`define LD4QHSP_D_F_Q_F 0.1
`define LD4QHSP_D_R_Q_R 0.1
`define LD4QHSP_D_GN_HOLD_posedge_posedge 0.1
`define LD4QHSP_D_GN_HOLD_negedge_posedge 0.1
`define LD4QHSP_D_GN_SETUP_posedge_posedge 0.1
`define LD4QHSP_D_GN_SETUP_negedge_posedge 0.1
`define LD4QHSP_GN_PWL 0.1
`define LD4QHSP_CD_PWL 0.1
`define LD4QHSP_CD_GN_REC_posedge_posedge 0.1
`define LD4QHSP_CD_GN_REM_posedge_posedge 0.1

module LD4QHSP (Q, D, GN, CD);

   output Q;
   input D;
   input GN;
   input CD;


   reg Notifier;


   U_LD_N_RN_NOTI u0 (IQ, D, GN, CD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if (!GN && CD) (D +=> Q) = (`LD4QHSP_D_R_Q_R,`LD4QHSP_D_F_Q_F);
      if(CD) (negedge GN => (Q +: D)) = (`LD4QHSP_GN_F_Q_R, `LD4QHSP_GN_F_Q_F);
      if(D && !GN) (posedge CD => (Q +: 1'b1)) = (`LD4QHSP_CD_R_Q_R,`LD4QHSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD4QHSP_CD_R_Q_R,`LD4QHSP_CD_F_Q_F);

	$setuphold(posedge GN &&& CD, posedge D, `LD4QHSP_D_GN_SETUP_posedge_posedge, `LD4QHSP_D_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& CD, negedge D, `LD4QHSP_D_GN_SETUP_negedge_posedge, `LD4QHSP_D_GN_HOLD_negedge_posedge, Notifier);

      $width(negedge GN, `LD4QHSP_GN_PWL, 0, Notifier);
      $width(negedge CD, `LD4QHSP_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge GN &&& D, `LD4QHSP_CD_GN_REC_posedge_posedge, Notifier);

	$hold(posedge GN &&& D, posedge CD, `LD4QHSP_CD_GN_REM_posedge_posedge, Notifier);

`else

      (D +=> Q) = (`LD4QHSP_D_R_Q_R,`LD4QHSP_D_F_Q_F);
      (negedge GN => (Q +: D)) = (`LD4QHSP_GN_F_Q_R, `LD4QHSP_GN_F_Q_F);
      (posedge CD => (Q +: 1'b1)) = (`LD4QHSP_CD_R_Q_R,`LD4QHSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD4QHSP_CD_R_Q_R,`LD4QHSP_CD_F_Q_F);
 
        $setuphold(posedge GN &&& CD, posedge D, `LD4QHSP_D_GN_SETUP_posedge_posedge, `LD4QHSP_D_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& CD, negedge D, `LD4QHSP_D_GN_SETUP_negedge_posedge, `LD4QHSP_D_GN_HOLD_negedge_posedge, Notifier);
 
      $width(negedge GN, `LD4QHSP_GN_PWL, 0, Notifier);
      $width(negedge CD, `LD4QHSP_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge GN &&& D, `LD4QHSP_CD_GN_REC_posedge_posedge, Notifier);
 
        $hold(posedge GN &&& D, posedge CD, `LD4QHSP_CD_GN_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD4QHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:17 and Version :1.1 //
 
//  START 
// CELL LD4QHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD4QHSX4_CD_F_Q_F 0.1
`define LD4QHSX4_CD_R_Q_R 0.1
`define LD4QHSX4_GN_F_Q_R 0.1
`define LD4QHSX4_GN_F_Q_F 0.1
`define LD4QHSX4_D_F_Q_F 0.1
`define LD4QHSX4_D_R_Q_R 0.1
`define LD4QHSX4_D_GN_HOLD_posedge_posedge 0.1
`define LD4QHSX4_D_GN_HOLD_negedge_posedge 0.1
`define LD4QHSX4_D_GN_SETUP_posedge_posedge 0.1
`define LD4QHSX4_D_GN_SETUP_negedge_posedge 0.1
`define LD4QHSX4_GN_PWL 0.1
`define LD4QHSX4_CD_PWL 0.1
`define LD4QHSX4_CD_GN_REC_posedge_posedge 0.1
`define LD4QHSX4_CD_GN_REM_posedge_posedge 0.1

module LD4QHSX4 (Q, D, GN, CD);

   output Q;
   input D;
   input GN;
   input CD;


   reg Notifier;


   U_LD_N_RN_NOTI u0 (IQ, D, GN, CD, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if (!GN && CD) (D +=> Q) = (`LD4QHSX4_D_R_Q_R,`LD4QHSX4_D_F_Q_F);
      if(CD) (negedge GN => (Q +: D)) = (`LD4QHSX4_GN_F_Q_R, `LD4QHSX4_GN_F_Q_F);
      if(D && !GN) (posedge CD => (Q +: 1'b1)) = (`LD4QHSX4_CD_R_Q_R,`LD4QHSX4_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD4QHSX4_CD_R_Q_R,`LD4QHSX4_CD_F_Q_F);

	$setuphold(posedge GN &&& CD, posedge D, `LD4QHSX4_D_GN_SETUP_posedge_posedge, `LD4QHSX4_D_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& CD, negedge D, `LD4QHSX4_D_GN_SETUP_negedge_posedge, `LD4QHSX4_D_GN_HOLD_negedge_posedge, Notifier);

      $width(negedge GN, `LD4QHSX4_GN_PWL, 0, Notifier);
      $width(negedge CD, `LD4QHSX4_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge GN &&& D, `LD4QHSX4_CD_GN_REC_posedge_posedge, Notifier);

	$hold(posedge GN &&& D, posedge CD, `LD4QHSX4_CD_GN_REM_posedge_posedge, Notifier);

`else

      (D +=> Q) = (`LD4QHSX4_D_R_Q_R,`LD4QHSX4_D_F_Q_F);
      (negedge GN => (Q +: D)) = (`LD4QHSX4_GN_F_Q_R, `LD4QHSX4_GN_F_Q_F);
      (posedge CD => (Q +: 1'b1)) = (`LD4QHSX4_CD_R_Q_R,`LD4QHSX4_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD4QHSX4_CD_R_Q_R,`LD4QHSX4_CD_F_Q_F);
 
        $setuphold(posedge GN &&& CD, posedge D, `LD4QHSX4_D_GN_SETUP_posedge_posedge, `LD4QHSX4_D_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& CD, negedge D, `LD4QHSX4_D_GN_SETUP_negedge_posedge, `LD4QHSX4_D_GN_HOLD_negedge_posedge, Notifier);
 
      $width(negedge GN, `LD4QHSX4_GN_PWL, 0, Notifier);
      $width(negedge CD, `LD4QHSX4_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge GN &&& D, `LD4QHSX4_CD_GN_REC_posedge_posedge, Notifier);
 
        $hold(posedge GN &&& D, posedge CD, `LD4QHSX4_CD_GN_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD4QHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:17 and Version :1.1 //
 
//  START 
// CELL LD4SHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD4SHS_TE_F_QN_R 0.1
`define LD4SHS_TE_R_QN_F 0.1
`define LD4SHS_TE_F_QN_F 0.1
`define LD4SHS_TE_R_QN_R 0.1
`define LD4SHS_TI_F_QN_R 0.1
`define LD4SHS_TI_R_QN_F 0.1
`define LD4SHS_CD_F_QN_R 0.1
`define LD4SHS_CD_R_QN_F 0.1
`define LD4SHS_GN_F_QN_F 0.1
`define LD4SHS_GN_F_QN_R 0.1
`define LD4SHS_D_F_QN_R 0.1
`define LD4SHS_D_R_QN_F 0.1
`define LD4SHS_TE_F_Q_F 0.1
`define LD4SHS_TE_R_Q_R 0.1
`define LD4SHS_TE_F_Q_R 0.1
`define LD4SHS_TE_R_Q_F 0.1
`define LD4SHS_TI_F_Q_F 0.1
`define LD4SHS_TI_R_Q_R 0.1
`define LD4SHS_CD_F_Q_F 0.1
`define LD4SHS_CD_R_Q_R 0.1
`define LD4SHS_GN_F_Q_R 0.1
`define LD4SHS_GN_F_Q_F 0.1
`define LD4SHS_D_F_Q_F 0.1
`define LD4SHS_D_R_Q_R 0.1
`define LD4SHS_CD_GN_REM_posedge_posedge 0.1
`define LD4SHS_CD_GN_REC_posedge_posedge 0.1
`define LD4SHS_CD_PWL 0.1
`define LD4SHS_GN_PWL 0.1
`define LD4SHS_D_GN_SETUP_posedge_posedge 0.1
`define LD4SHS_D_GN_SETUP_negedge_posedge 0.1
`define LD4SHS_D_GN_HOLD_posedge_posedge 0.1
`define LD4SHS_D_GN_HOLD_negedge_posedge 0.1
`define LD4SHS_TI_GN_SETUP_posedge_posedge 0.1
`define LD4SHS_TI_GN_SETUP_negedge_posedge 0.1
`define LD4SHS_TI_GN_HOLD_posedge_posedge 0.1
`define LD4SHS_TI_GN_HOLD_negedge_posedge 0.1
`define LD4SHS_TE_GN_SETUP_posedge_posedge 0.1
`define LD4SHS_TE_GN_SETUP_negedge_posedge 0.1
`define LD4SHS_TE_GN_HOLD_posedge_posedge 0.1
`define LD4SHS_TE_GN_HOLD_negedge_posedge 0.1

module LD4SHS (Q, QN, D, GN, CD, TI, TE);

   output Q;
   output QN;
   input D;
   input GN;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_LD_N_RN_NOTI u1 (   // Verilog Seq UDP
      IQ, Mux21DTITE_, GN, CD, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);



`ifdef functional
`else
   not  (TEX, TE);
   and  (AndCDTEX_, CD, TEX);
   and  (AndCDTE_, CD, TE);
   xor  (XorDTI_, D, TI);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   specify
`ifdef verifault

      if (!D && !GN && TI) (TE -=> QN) = (`LD4SHS_TE_F_QN_R,`LD4SHS_TE_R_QN_F);
      if (D && !GN && !TI) (TE +=> QN) = (`LD4SHS_TE_R_QN_R,`LD4SHS_TE_F_QN_F);
      if (!GN && CD && TE) (TI -=> QN) = (`LD4SHS_TI_F_QN_R,`LD4SHS_TI_R_QN_F);
      if (!GN && CD && !TE) (D -=> QN) = (`LD4SHS_D_F_QN_R,`LD4SHS_D_R_QN_F);
      if (!D && !GN && TI) (TE +=> Q) = (`LD4SHS_TE_R_Q_R,`LD4SHS_TE_F_Q_F);
      if (D && !GN && !TI) (TE -=> Q) = (`LD4SHS_TE_F_Q_R,`LD4SHS_TE_R_Q_F);
      if (!GN && CD && TE) (TI +=> Q) = (`LD4SHS_TI_R_Q_R,`LD4SHS_TI_F_Q_F);
      if (!GN && CD && !TE) (D +=> Q) = (`LD4SHS_D_R_Q_R,`LD4SHS_D_F_Q_F);
      if(!TE) (negedge GN => (Q +: D)) = (`LD4SHS_GN_F_Q_R, `LD4SHS_GN_F_Q_F);
      if(TE) (negedge GN => (Q +: TI)) = (`LD4SHS_GN_F_Q_R, `LD4SHS_GN_F_Q_F);
      if(!D && TI) (negedge GN => (Q +: TE)) = (`LD4SHS_GN_F_Q_R, `LD4SHS_GN_F_Q_F);
      if(!TI && D) (negedge GN => (Q -: TE)) = (`LD4SHS_GN_F_Q_R, `LD4SHS_GN_F_Q_F);
      if(!TE) (negedge GN => (QN -: D)) = (`LD4SHS_GN_F_QN_R, `LD4SHS_GN_F_QN_F);
      if(TE) (negedge GN => (QN -: TI)) = (`LD4SHS_GN_F_QN_R, `LD4SHS_GN_F_QN_F);
      if(!D && TI) (negedge GN => (QN -: TE)) = (`LD4SHS_GN_F_QN_R, `LD4SHS_GN_F_QN_F);
      if(!TI && D) (negedge GN => (QN +: TE)) = (`LD4SHS_GN_F_QN_R, `LD4SHS_GN_F_QN_F);
      if(D && !GN && !TE || !GN && TI && TE) (posedge CD => (Q +: 1'b1)) = (`LD4SHS_CD_R_Q_R,`LD4SHS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD4SHS_CD_R_Q_R,`LD4SHS_CD_F_Q_F);
      if(D && !GN && !TE || !GN && TI && TE) (posedge CD => (QN +: 1'b0)) = (`LD4SHS_CD_F_QN_R,`LD4SHS_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`LD4SHS_CD_F_QN_R,`LD4SHS_CD_R_QN_F);

	$setuphold(posedge GN &&& AndXorDTI_CD_, posedge TE, `LD4SHS_TE_GN_SETUP_posedge_posedge, `LD4SHS_TE_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& AndXorDTI_CD_, negedge TE, `LD4SHS_TE_GN_SETUP_negedge_posedge, `LD4SHS_TE_GN_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge GN &&& AndCDTE_, posedge TI, `LD4SHS_TI_GN_SETUP_posedge_posedge, `LD4SHS_TI_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& AndCDTE_, negedge TI, `LD4SHS_TI_GN_SETUP_negedge_posedge, `LD4SHS_TI_GN_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge GN &&& AndCDTEX_, posedge D, `LD4SHS_D_GN_SETUP_posedge_posedge, `LD4SHS_D_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& AndCDTEX_, negedge D, `LD4SHS_D_GN_SETUP_negedge_posedge, `LD4SHS_D_GN_HOLD_negedge_posedge, Notifier);

      $width(negedge GN, `LD4SHS_GN_PWL, 0, Notifier);
      $width(negedge CD, `LD4SHS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge GN &&& Mux21DTITE_, `LD4SHS_CD_GN_REC_posedge_posedge, Notifier);

	$hold(posedge GN &&& Mux21DTITE_, posedge CD, `LD4SHS_CD_GN_REM_posedge_posedge, Notifier);

`else
      if (!D && !GN && TI) (TE -=> QN) = (`LD4SHS_TE_F_QN_R,`LD4SHS_TE_R_QN_F);
      if (D && !GN && !TI) (TE +=> QN) = (`LD4SHS_TE_R_QN_R,`LD4SHS_TE_F_QN_F);
       (TI -=> QN) = (`LD4SHS_TI_F_QN_R,`LD4SHS_TI_R_QN_F);
       (D -=> QN) = (`LD4SHS_D_F_QN_R,`LD4SHS_D_R_QN_F);
      if (!D && !GN && TI) (TE +=> Q) = (`LD4SHS_TE_R_Q_R,`LD4SHS_TE_F_Q_F);
      if (D && !GN && !TI) (TE -=> Q) = (`LD4SHS_TE_F_Q_R,`LD4SHS_TE_R_Q_F);
      (TI +=> Q) = (`LD4SHS_TI_R_Q_R,`LD4SHS_TI_F_Q_F);
      (D +=> Q) = (`LD4SHS_D_R_Q_R,`LD4SHS_D_F_Q_F);
      (negedge GN => (Q +: Mux21DTITE_)) = (`LD4SHS_GN_F_Q_R, `LD4SHS_GN_F_Q_F);
      (negedge GN => (QN -: Mux21DTITE_)) = (`LD4SHS_GN_F_QN_R, `LD4SHS_GN_F_QN_F);
      (posedge CD => (Q +: 1'b1)) = (`LD4SHS_CD_R_Q_R,`LD4SHS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD4SHS_CD_R_Q_R,`LD4SHS_CD_F_Q_F);
      (posedge CD => (QN +: 1'b0)) = (`LD4SHS_CD_F_QN_R,`LD4SHS_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`LD4SHS_CD_F_QN_R,`LD4SHS_CD_R_QN_F);
 
        $setuphold(posedge GN &&& AndXorDTI_CD_, posedge TE, `LD4SHS_TE_GN_SETUP_posedge_posedge, `LD4SHS_TE_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& AndXorDTI_CD_, negedge TE, `LD4SHS_TE_GN_SETUP_negedge_posedge, `LD4SHS_TE_GN_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge GN &&& AndCDTE_, posedge TI, `LD4SHS_TI_GN_SETUP_posedge_posedge, `LD4SHS_TI_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& AndCDTE_, negedge TI, `LD4SHS_TI_GN_SETUP_negedge_posedge, `LD4SHS_TI_GN_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge GN &&& AndCDTEX_, posedge D, `LD4SHS_D_GN_SETUP_posedge_posedge, `LD4SHS_D_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& AndCDTEX_, negedge D, `LD4SHS_D_GN_SETUP_negedge_posedge, `LD4SHS_D_GN_HOLD_negedge_posedge, Notifier);
 
      $width(negedge GN, `LD4SHS_GN_PWL, 0, Notifier);
      $width(negedge CD, `LD4SHS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge GN &&& Mux21DTITE_, `LD4SHS_CD_GN_REC_posedge_posedge, Notifier);
 
        $hold(posedge GN &&& Mux21DTITE_, posedge CD, `LD4SHS_CD_GN_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD4SHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:23 and Version :1.1 //
 
//  START 
// CELL LD4SQHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD4SQHS_TE_F_Q_F 0.1
`define LD4SQHS_TE_R_Q_R 0.1
`define LD4SQHS_TE_F_Q_R 0.1
`define LD4SQHS_TE_R_Q_F 0.1
`define LD4SQHS_TI_F_Q_F 0.1
`define LD4SQHS_TI_R_Q_R 0.1
`define LD4SQHS_CD_F_Q_F 0.1
`define LD4SQHS_CD_R_Q_R 0.1
`define LD4SQHS_GN_F_Q_R 0.1
`define LD4SQHS_GN_F_Q_F 0.1
`define LD4SQHS_D_F_Q_F 0.1
`define LD4SQHS_D_R_Q_R 0.1
`define LD4SQHS_TE_GN_HOLD_posedge_posedge 0.1
`define LD4SQHS_TE_GN_HOLD_negedge_posedge 0.1
`define LD4SQHS_TE_GN_SETUP_posedge_posedge 0.1
`define LD4SQHS_TE_GN_SETUP_negedge_posedge 0.1
`define LD4SQHS_TI_GN_HOLD_posedge_posedge 0.1
`define LD4SQHS_TI_GN_HOLD_negedge_posedge 0.1
`define LD4SQHS_TI_GN_SETUP_posedge_posedge 0.1
`define LD4SQHS_TI_GN_SETUP_negedge_posedge 0.1
`define LD4SQHS_D_GN_HOLD_posedge_posedge 0.1
`define LD4SQHS_D_GN_HOLD_negedge_posedge 0.1
`define LD4SQHS_D_GN_SETUP_posedge_posedge 0.1
`define LD4SQHS_D_GN_SETUP_negedge_posedge 0.1
`define LD4SQHS_GN_PWL 0.1
`define LD4SQHS_CD_PWL 0.1
`define LD4SQHS_CD_GN_REC_posedge_posedge 0.1
`define LD4SQHS_CD_GN_REM_posedge_posedge 0.1

module LD4SQHS (Q, D, GN, CD, TI, TE);

   output Q;
   input D;
   input GN;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_LD_N_RN_NOTI u1 (IQ, Mux21DTITE_, GN, CD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if (!D && !GN && TI) (TE +=> Q) = (`LD4SQHS_TE_R_Q_R,`LD4SQHS_TE_F_Q_F);
      if (D && !GN && !TI) (TE -=> Q) = (`LD4SQHS_TE_F_Q_R,`LD4SQHS_TE_R_Q_F);
      if (!GN && CD && TE) (TI +=> Q) = (`LD4SQHS_TI_R_Q_R,`LD4SQHS_TI_F_Q_F);
      if (!GN && CD && !TE) (D +=> Q) = (`LD4SQHS_D_R_Q_R,`LD4SQHS_D_F_Q_F);
      if(!TE && CD) (negedge GN => (Q +: D)) = (`LD4SQHS_GN_F_Q_R, `LD4SQHS_GN_F_Q_F);
      if(TE && CD) (negedge GN => (Q +: TI)) = (`LD4SQHS_GN_F_Q_R, `LD4SQHS_GN_F_Q_F);
      if(!D && TI && CD) (negedge GN => (Q +: TE)) = (`LD4SQHS_GN_F_Q_R, `LD4SQHS_GN_F_Q_F);
      if(!TI && D && CD) (negedge GN => (Q -: TE)) = (`LD4SQHS_GN_F_Q_R, `LD4SQHS_GN_F_Q_F);
      if(D && !GN && !TE || !GN && TI && TE) (posedge CD => (Q +: 1'b1)) = (`LD4SQHS_CD_R_Q_R,`LD4SQHS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD4SQHS_CD_R_Q_R,`LD4SQHS_CD_F_Q_F);

	$setuphold(posedge GN &&& AndXorDTI_CD_, posedge TE, `LD4SQHS_TE_GN_SETUP_posedge_posedge, `LD4SQHS_TE_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& AndXorDTI_CD_, negedge TE, `LD4SQHS_TE_GN_SETUP_negedge_posedge, `LD4SQHS_TE_GN_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge GN &&& AndCDTE_, posedge TI, `LD4SQHS_TI_GN_SETUP_posedge_posedge, `LD4SQHS_TI_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& AndCDTE_, negedge TI, `LD4SQHS_TI_GN_SETUP_negedge_posedge, `LD4SQHS_TI_GN_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge GN &&& AndCDTEX_, posedge D, `LD4SQHS_D_GN_SETUP_posedge_posedge, `LD4SQHS_D_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& AndCDTEX_, negedge D, `LD4SQHS_D_GN_SETUP_negedge_posedge, `LD4SQHS_D_GN_HOLD_negedge_posedge, Notifier);

      $width(negedge GN, `LD4SQHS_GN_PWL, 0, Notifier);
      $width(negedge CD, `LD4SQHS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge GN &&& Mux21DTITE_, `LD4SQHS_CD_GN_REC_posedge_posedge, Notifier);

	$hold(posedge GN &&& Mux21DTITE_, posedge CD, `LD4SQHS_CD_GN_REM_posedge_posedge, Notifier);

`else

     if (!D && !GN && TI) (TE +=>Q) = (`LD4SQHS_TE_R_Q_R,`LD4SQHS_TE_F_Q_F);
      if (D && !GN && !TI) (TE -=> Q) = (`LD4SQHS_TE_F_Q_R,`LD4SQHS_TE_R_Q_F);
      (TI +=>Q ) = (`LD4SQHS_TI_R_Q_R,`LD4SQHS_TI_F_Q_F);
      (D +=> Q) = (`LD4SQHS_D_R_Q_R,`LD4SQHS_D_F_Q_F);
      (negedge GN => (Q +: Mux21DTITE_)) = (`LD4SQHS_GN_F_Q_R, `LD4SQHS_GN_F_Q_F);
      (posedge CD => (Q +: 1'b1)) = (`LD4SQHS_CD_R_Q_R,`LD4SQHS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD4SQHS_CD_R_Q_R,`LD4SQHS_CD_F_Q_F);
 
        $setuphold(posedge GN &&& AndXorDTI_CD_, posedge TE, `LD4SQHS_TE_GN_SETUP_posedge_posedge, `LD4SQHS_TE_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& AndXorDTI_CD_, negedge TE, `LD4SQHS_TE_GN_SETUP_negedge_posedge, `LD4SQHS_TE_GN_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge GN &&& AndCDTE_, posedge TI, `LD4SQHS_TI_GN_SETUP_posedge_posedge, `LD4SQHS_TI_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& AndCDTE_, negedge TI, `LD4SQHS_TI_GN_SETUP_negedge_posedge, `LD4SQHS_TI_GN_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge GN &&& AndCDTEX_, posedge D, `LD4SQHS_D_GN_SETUP_posedge_posedge, `LD4SQHS_D_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& AndCDTEX_, negedge D, `LD4SQHS_D_GN_SETUP_negedge_posedge, `LD4SQHS_D_GN_HOLD_negedge_posedge, Notifier);
 
      $width(negedge GN, `LD4SQHS_GN_PWL, 0, Notifier);
      $width(negedge CD, `LD4SQHS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge GN &&& Mux21DTITE_, `LD4SQHS_CD_GN_REC_posedge_posedge, Notifier);
 
        $hold(posedge GN &&& Mux21DTITE_, posedge CD, `LD4SQHS_CD_GN_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD4SQHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:23 and Version :1.1 //
 
//  START 
// CELL LD4SQHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD4SQHSP_TE_F_Q_F 0.1
`define LD4SQHSP_TE_R_Q_R 0.1
`define LD4SQHSP_TE_F_Q_R 0.1
`define LD4SQHSP_TE_R_Q_F 0.1
`define LD4SQHSP_TI_F_Q_F 0.1
`define LD4SQHSP_TI_R_Q_R 0.1
`define LD4SQHSP_CD_F_Q_F 0.1
`define LD4SQHSP_CD_R_Q_R 0.1
`define LD4SQHSP_GN_F_Q_R 0.1
`define LD4SQHSP_GN_F_Q_F 0.1
`define LD4SQHSP_D_F_Q_F 0.1
`define LD4SQHSP_D_R_Q_R 0.1
`define LD4SQHSP_TE_GN_HOLD_posedge_posedge 0.1
`define LD4SQHSP_TE_GN_HOLD_negedge_posedge 0.1
`define LD4SQHSP_TE_GN_SETUP_posedge_posedge 0.1
`define LD4SQHSP_TE_GN_SETUP_negedge_posedge 0.1
`define LD4SQHSP_TI_GN_HOLD_posedge_posedge 0.1
`define LD4SQHSP_TI_GN_HOLD_negedge_posedge 0.1
`define LD4SQHSP_TI_GN_SETUP_posedge_posedge 0.1
`define LD4SQHSP_TI_GN_SETUP_negedge_posedge 0.1
`define LD4SQHSP_D_GN_HOLD_posedge_posedge 0.1
`define LD4SQHSP_D_GN_HOLD_negedge_posedge 0.1
`define LD4SQHSP_D_GN_SETUP_posedge_posedge 0.1
`define LD4SQHSP_D_GN_SETUP_negedge_posedge 0.1
`define LD4SQHSP_GN_PWL 0.1
`define LD4SQHSP_CD_PWL 0.1
`define LD4SQHSP_CD_GN_REC_posedge_posedge 0.1
`define LD4SQHSP_CD_GN_REM_posedge_posedge 0.1

module LD4SQHSP (Q, D, GN, CD, TI, TE);

   output Q;
   input D;
   input GN;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_LD_N_RN_NOTI u1 (IQ, Mux21DTITE_, GN, CD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if (!D && !GN && TI) (TE +=> Q) = (`LD4SQHSP_TE_R_Q_R,`LD4SQHSP_TE_F_Q_F);
      if (D && !GN && !TI) (TE -=> Q) = (`LD4SQHSP_TE_F_Q_R,`LD4SQHSP_TE_R_Q_F);
      if (!GN && CD && TE) (TI +=> Q) = (`LD4SQHSP_TI_R_Q_R,`LD4SQHSP_TI_F_Q_F);
      if (!GN && CD && !TE) (D +=> Q) = (`LD4SQHSP_D_R_Q_R,`LD4SQHSP_D_F_Q_F);
      if(!TE && CD) (negedge GN => (Q +: D)) = (`LD4SQHSP_GN_F_Q_R, `LD4SQHSP_GN_F_Q_F);
      if(TE && CD) (negedge GN => (Q +: TI)) = (`LD4SQHSP_GN_F_Q_R, `LD4SQHSP_GN_F_Q_F);
      if(!D && TI && CD) (negedge GN => (Q +: TE)) = (`LD4SQHSP_GN_F_Q_R, `LD4SQHSP_GN_F_Q_F);
      if(!TI && D && CD) (negedge GN => (Q -: TE)) = (`LD4SQHSP_GN_F_Q_R, `LD4SQHSP_GN_F_Q_F);
      if(D && !GN && !TE || !GN && TI && TE) (posedge CD => (Q +: 1'b1)) = (`LD4SQHSP_CD_R_Q_R,`LD4SQHSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD4SQHSP_CD_R_Q_R,`LD4SQHSP_CD_F_Q_F);

	$setuphold(posedge GN &&& AndXorDTI_CD_, posedge TE, `LD4SQHSP_TE_GN_SETUP_posedge_posedge, `LD4SQHSP_TE_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& AndXorDTI_CD_, negedge TE, `LD4SQHSP_TE_GN_SETUP_negedge_posedge, `LD4SQHSP_TE_GN_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge GN &&& AndCDTE_, posedge TI, `LD4SQHSP_TI_GN_SETUP_posedge_posedge, `LD4SQHSP_TI_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& AndCDTE_, negedge TI, `LD4SQHSP_TI_GN_SETUP_negedge_posedge, `LD4SQHSP_TI_GN_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge GN &&& AndCDTEX_, posedge D, `LD4SQHSP_D_GN_SETUP_posedge_posedge, `LD4SQHSP_D_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& AndCDTEX_, negedge D, `LD4SQHSP_D_GN_SETUP_negedge_posedge, `LD4SQHSP_D_GN_HOLD_negedge_posedge, Notifier);

      $width(negedge GN, `LD4SQHSP_GN_PWL, 0, Notifier);
      $width(negedge CD, `LD4SQHSP_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge GN &&& Mux21DTITE_, `LD4SQHSP_CD_GN_REC_posedge_posedge, Notifier);

	$hold(posedge GN &&& Mux21DTITE_, posedge CD, `LD4SQHSP_CD_GN_REM_posedge_posedge, Notifier);

`else

     if (!D && !GN && TI) (TE +=>Q) = (`LD4SQHSP_TE_R_Q_R,`LD4SQHSP_TE_F_Q_F);
      if (D && !GN && !TI) (TE -=> Q) = (`LD4SQHSP_TE_F_Q_R,`LD4SQHSP_TE_R_Q_F);
      (TI +=>Q ) = (`LD4SQHSP_TI_R_Q_R,`LD4SQHSP_TI_F_Q_F);
      (D +=> Q) = (`LD4SQHSP_D_R_Q_R,`LD4SQHSP_D_F_Q_F);
      (negedge GN => (Q +: Mux21DTITE_)) = (`LD4SQHSP_GN_F_Q_R, `LD4SQHSP_GN_F_Q_F);
      (posedge CD => (Q +: 1'b1)) = (`LD4SQHSP_CD_R_Q_R,`LD4SQHSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD4SQHSP_CD_R_Q_R,`LD4SQHSP_CD_F_Q_F);
 
        $setuphold(posedge GN &&& AndXorDTI_CD_, posedge TE, `LD4SQHSP_TE_GN_SETUP_posedge_posedge, `LD4SQHSP_TE_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& AndXorDTI_CD_, negedge TE, `LD4SQHSP_TE_GN_SETUP_negedge_posedge, `LD4SQHSP_TE_GN_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge GN &&& AndCDTE_, posedge TI, `LD4SQHSP_TI_GN_SETUP_posedge_posedge, `LD4SQHSP_TI_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& AndCDTE_, negedge TI, `LD4SQHSP_TI_GN_SETUP_negedge_posedge, `LD4SQHSP_TI_GN_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge GN &&& AndCDTEX_, posedge D, `LD4SQHSP_D_GN_SETUP_posedge_posedge, `LD4SQHSP_D_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& AndCDTEX_, negedge D, `LD4SQHSP_D_GN_SETUP_negedge_posedge, `LD4SQHSP_D_GN_HOLD_negedge_posedge, Notifier);
 
      $width(negedge GN, `LD4SQHSP_GN_PWL, 0, Notifier);
      $width(negedge CD, `LD4SQHSP_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge GN &&& Mux21DTITE_, `LD4SQHSP_CD_GN_REC_posedge_posedge, Notifier);
 
        $hold(posedge GN &&& Mux21DTITE_, posedge CD, `LD4SQHSP_CD_GN_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD4SQHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:23 and Version :1.1 //
 
//  START 
// CELL LD4SQHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD4SQHSX4_TE_F_Q_F 0.1
`define LD4SQHSX4_TE_R_Q_R 0.1
`define LD4SQHSX4_TE_F_Q_R 0.1
`define LD4SQHSX4_TE_R_Q_F 0.1
`define LD4SQHSX4_TI_F_Q_F 0.1
`define LD4SQHSX4_TI_R_Q_R 0.1
`define LD4SQHSX4_CD_F_Q_F 0.1
`define LD4SQHSX4_CD_R_Q_R 0.1
`define LD4SQHSX4_GN_F_Q_R 0.1
`define LD4SQHSX4_GN_F_Q_F 0.1
`define LD4SQHSX4_D_F_Q_F 0.1
`define LD4SQHSX4_D_R_Q_R 0.1
`define LD4SQHSX4_TE_GN_HOLD_posedge_posedge 0.1
`define LD4SQHSX4_TE_GN_HOLD_negedge_posedge 0.1
`define LD4SQHSX4_TE_GN_SETUP_posedge_posedge 0.1
`define LD4SQHSX4_TE_GN_SETUP_negedge_posedge 0.1
`define LD4SQHSX4_TI_GN_HOLD_posedge_posedge 0.1
`define LD4SQHSX4_TI_GN_HOLD_negedge_posedge 0.1
`define LD4SQHSX4_TI_GN_SETUP_posedge_posedge 0.1
`define LD4SQHSX4_TI_GN_SETUP_negedge_posedge 0.1
`define LD4SQHSX4_D_GN_HOLD_posedge_posedge 0.1
`define LD4SQHSX4_D_GN_HOLD_negedge_posedge 0.1
`define LD4SQHSX4_D_GN_SETUP_posedge_posedge 0.1
`define LD4SQHSX4_D_GN_SETUP_negedge_posedge 0.1
`define LD4SQHSX4_GN_PWL 0.1
`define LD4SQHSX4_CD_PWL 0.1
`define LD4SQHSX4_CD_GN_REC_posedge_posedge 0.1
`define LD4SQHSX4_CD_GN_REM_posedge_posedge 0.1

module LD4SQHSX4 (Q, D, GN, CD, TI, TE);

   output Q;
   input D;
   input GN;
   input CD;
   input TI;
   input TE;


   reg Notifier;

   U_MUX2  u0 (Mux21DTITE_, D, TI, TE);

   U_LD_N_RN_NOTI u1 (IQ, Mux21DTITE_, GN, CD, Notifier);

   buf  u2 (Q, IQ);



`ifdef functional
`else
   and  (AndCDTEX_, CD, TEX);
   not  (TEX, TE);
   and  (AndCDTE_, CD, TE);
   and  (AndXorDTI_CD_, XorDTI_, CD);
   xor  (XorDTI_, D, TI);
   // if(TE==0) DorTIonTE = D; else DorTIonTE = TI ;
   and  (AndTETI, TE, TI);
   and  (AndTEXD, TEX, D);
   or   (DorTIonTE, AndTETI, AndTEXD);

   specify
`ifdef verifault

      if (!D && !GN && TI) (TE +=> Q) = (`LD4SQHSX4_TE_R_Q_R,`LD4SQHSX4_TE_F_Q_F);
      if (D && !GN && !TI) (TE -=> Q) = (`LD4SQHSX4_TE_F_Q_R,`LD4SQHSX4_TE_R_Q_F);
      if (!GN && CD && TE) (TI +=> Q) = (`LD4SQHSX4_TI_R_Q_R,`LD4SQHSX4_TI_F_Q_F);
      if (!GN && CD && !TE) (D +=> Q) = (`LD4SQHSX4_D_R_Q_R,`LD4SQHSX4_D_F_Q_F);
      if(!TE && CD) (negedge GN => (Q +: D)) = (`LD4SQHSX4_GN_F_Q_R, `LD4SQHSX4_GN_F_Q_F);
      if(TE && CD) (negedge GN => (Q +: TI)) = (`LD4SQHSX4_GN_F_Q_R, `LD4SQHSX4_GN_F_Q_F);
      if(!D && TI && CD) (negedge GN => (Q +: TE)) = (`LD4SQHSX4_GN_F_Q_R, `LD4SQHSX4_GN_F_Q_F);
      if(!TI && D && CD) (negedge GN => (Q -: TE)) = (`LD4SQHSX4_GN_F_Q_R, `LD4SQHSX4_GN_F_Q_F);
      if(D && !GN && !TE || !GN && TI && TE) (posedge CD => (Q +: 1'b1)) = (`LD4SQHSX4_CD_R_Q_R,`LD4SQHSX4_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD4SQHSX4_CD_R_Q_R,`LD4SQHSX4_CD_F_Q_F);

	$setuphold(posedge GN &&& AndXorDTI_CD_, posedge TE, `LD4SQHSX4_TE_GN_SETUP_posedge_posedge, `LD4SQHSX4_TE_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& AndXorDTI_CD_, negedge TE, `LD4SQHSX4_TE_GN_SETUP_negedge_posedge, `LD4SQHSX4_TE_GN_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge GN &&& AndCDTE_, posedge TI, `LD4SQHSX4_TI_GN_SETUP_posedge_posedge, `LD4SQHSX4_TI_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& AndCDTE_, negedge TI, `LD4SQHSX4_TI_GN_SETUP_negedge_posedge, `LD4SQHSX4_TI_GN_HOLD_negedge_posedge, Notifier);

	$setuphold(posedge GN &&& AndCDTEX_, posedge D, `LD4SQHSX4_D_GN_SETUP_posedge_posedge, `LD4SQHSX4_D_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& AndCDTEX_, negedge D, `LD4SQHSX4_D_GN_SETUP_negedge_posedge, `LD4SQHSX4_D_GN_HOLD_negedge_posedge, Notifier);

      $width(negedge GN, `LD4SQHSX4_GN_PWL, 0, Notifier);
      $width(negedge CD, `LD4SQHSX4_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge GN &&& Mux21DTITE_, `LD4SQHSX4_CD_GN_REC_posedge_posedge, Notifier);

	$hold(posedge GN &&& Mux21DTITE_, posedge CD, `LD4SQHSX4_CD_GN_REM_posedge_posedge, Notifier);

`else

     if (!D && !GN && TI) (TE +=>Q) = (`LD4SQHSX4_TE_R_Q_R,`LD4SQHSX4_TE_F_Q_F);
      if (D && !GN && !TI) (TE -=> Q) = (`LD4SQHSX4_TE_F_Q_R,`LD4SQHSX4_TE_R_Q_F);
      (TI +=>Q ) = (`LD4SQHSX4_TI_R_Q_R,`LD4SQHSX4_TI_F_Q_F);
      (D +=> Q) = (`LD4SQHSX4_D_R_Q_R,`LD4SQHSX4_D_F_Q_F);
      (negedge GN => (Q +: Mux21DTITE_)) = (`LD4SQHSX4_GN_F_Q_R, `LD4SQHSX4_GN_F_Q_F);
      (posedge CD => (Q +: 1'b1)) = (`LD4SQHSX4_CD_R_Q_R,`LD4SQHSX4_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD4SQHSX4_CD_R_Q_R,`LD4SQHSX4_CD_F_Q_F);
 
        $setuphold(posedge GN &&& AndXorDTI_CD_, posedge TE, `LD4SQHSX4_TE_GN_SETUP_posedge_posedge, `LD4SQHSX4_TE_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& AndXorDTI_CD_, negedge TE, `LD4SQHSX4_TE_GN_SETUP_negedge_posedge, `LD4SQHSX4_TE_GN_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge GN &&& AndCDTE_, posedge TI, `LD4SQHSX4_TI_GN_SETUP_posedge_posedge, `LD4SQHSX4_TI_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& AndCDTE_, negedge TI, `LD4SQHSX4_TI_GN_SETUP_negedge_posedge, `LD4SQHSX4_TI_GN_HOLD_negedge_posedge, Notifier);
 
        $setuphold(posedge GN &&& AndCDTEX_, posedge D, `LD4SQHSX4_D_GN_SETUP_posedge_posedge, `LD4SQHSX4_D_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& AndCDTEX_, negedge D, `LD4SQHSX4_D_GN_SETUP_negedge_posedge, `LD4SQHSX4_D_GN_HOLD_negedge_posedge, Notifier);
 
      $width(negedge GN, `LD4SQHSX4_GN_PWL, 0, Notifier);
      $width(negedge CD, `LD4SQHSX4_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge GN &&& Mux21DTITE_, `LD4SQHSX4_CD_GN_REC_posedge_posedge, Notifier);
 
        $hold(posedge GN &&& Mux21DTITE_, posedge CD, `LD4SQHSX4_CD_GN_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD4SQHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:23 and Version :1.1 //
 
//  START 
// CELL LD5HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD5HS_SD_F_QN_F 0.1
`define LD5HS_SD_R_QN_R 0.1
`define LD5HS_G_R_QN_F 0.1
`define LD5HS_G_R_QN_R 0.1
`define LD5HS_D_F_QN_R 0.1
`define LD5HS_D_R_QN_F 0.1
`define LD5HS_SD_F_Q_R 0.1
`define LD5HS_SD_R_Q_F 0.1
`define LD5HS_G_R_Q_R 0.1
`define LD5HS_G_R_Q_F 0.1
`define LD5HS_D_F_Q_F 0.1
`define LD5HS_D_R_Q_R 0.1
`define LD5HS_D_G_HOLD_posedge_negedge 0.1
`define LD5HS_D_G_HOLD_negedge_negedge 0.1
`define LD5HS_D_G_SETUP_posedge_negedge 0.1
`define LD5HS_D_G_SETUP_negedge_negedge 0.1
`define LD5HS_G_PWH 0.1
`define LD5HS_SD_PWL 0.1
`define LD5HS_SD_G_REC_posedge_negedge 0.1
`define LD5HS_SD_G_REM_posedge_negedge 0.1

module LD5HS (Q, QN, D, G, SD);

   output Q;
   output QN;
   input D;
   input G;
   input SD;


   reg Notifier;


   U_LD_P_SN_NOTI u0 (IQ, D, G, SD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   not  (GX, G);
   not  (D_, D);
   specify
`ifdef verifault

      if (G && SD) (D -=> QN) = (`LD5HS_D_F_QN_R,`LD5HS_D_R_QN_F);
      if (G && SD) (D +=> Q) = (`LD5HS_D_R_Q_R,`LD5HS_D_F_Q_F);
      if(SD) (posedge G => (Q +: D)) = (`LD5HS_G_R_Q_R, `LD5HS_G_R_Q_F);
      if(SD) (posedge G => (QN -: D)) = (`LD5HS_G_R_QN_R, `LD5HS_G_R_QN_F);
      if(!D && G) (posedge SD => (Q +: 1'b0)) = (`LD5HS_SD_F_Q_R,`LD5HS_SD_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`LD5HS_SD_F_Q_R,`LD5HS_SD_R_Q_F);
      if(!D && G) (posedge SD => (QN +: 1'b1)) = (`LD5HS_SD_R_QN_R,`LD5HS_SD_F_QN_F);
      (negedge SD => (QN +: 1'b0)) = (`LD5HS_SD_R_QN_R,`LD5HS_SD_F_QN_F);

	$setuphold(negedge G &&& SD, posedge D, `LD5HS_D_G_SETUP_posedge_negedge, `LD5HS_D_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& SD, negedge D, `LD5HS_D_G_SETUP_negedge_negedge, `LD5HS_D_G_HOLD_negedge_negedge, Notifier);

      $width(posedge G, `LD5HS_G_PWH, 0, Notifier);
      $width(negedge SD, `LD5HS_SD_PWL, 0, Notifier);
	$recovery(posedge SD, negedge G &&& D_, `LD5HS_SD_G_REC_posedge_negedge, Notifier);

	$hold(negedge G &&& D_, posedge SD, `LD5HS_SD_G_REM_posedge_negedge, Notifier);
`else

      (D -=> QN) = (`LD5HS_D_F_QN_R,`LD5HS_D_R_QN_F);
      (D +=> Q) = (`LD5HS_D_R_Q_R,`LD5HS_D_F_Q_F);
      (posedge G => (Q +: D)) = (`LD5HS_G_R_Q_R, `LD5HS_G_R_Q_F);
            (posedge G => (QN -: D)) = (`LD5HS_G_R_QN_R, `LD5HS_G_R_QN_F);
      (posedge SD => (Q +: 1'b0)) = (`LD5HS_SD_F_Q_R,`LD5HS_SD_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`LD5HS_SD_F_Q_R,`LD5HS_SD_R_Q_F);
      (posedge SD => (QN +: 1'b1)) = (`LD5HS_SD_R_QN_R,`LD5HS_SD_F_QN_F);
      (negedge SD => (QN +: 1'b0)) = (`LD5HS_SD_R_QN_R,`LD5HS_SD_F_QN_F);
 
        $setuphold(negedge G &&& SD, posedge D, `LD5HS_D_G_SETUP_posedge_negedge, `LD5HS_D_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& SD, negedge D, `LD5HS_D_G_SETUP_negedge_negedge, `LD5HS_D_G_HOLD_negedge_negedge, Notifier);
 
      $width(posedge G, `LD5HS_G_PWH, 0, Notifier);
      $width(negedge SD, `LD5HS_SD_PWL, 0, Notifier);
        $recovery(posedge SD, negedge G &&& D_, `LD5HS_SD_G_REC_posedge_negedge, Notifier);
 
        $hold(negedge G &&& D_, posedge SD, `LD5HS_SD_G_REM_posedge_negedge, Notifier);

`endif
   endspecify
`endif


endmodule // LD5HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:27 and Version :1.1 //
 
//  START 
// CELL LD5HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD5HSP_SD_F_QN_F 0.1
`define LD5HSP_SD_R_QN_R 0.1
`define LD5HSP_G_R_QN_F 0.1
`define LD5HSP_G_R_QN_R 0.1
`define LD5HSP_D_F_QN_R 0.1
`define LD5HSP_D_R_QN_F 0.1
`define LD5HSP_SD_F_Q_R 0.1
`define LD5HSP_SD_R_Q_F 0.1
`define LD5HSP_G_R_Q_R 0.1
`define LD5HSP_G_R_Q_F 0.1
`define LD5HSP_D_F_Q_F 0.1
`define LD5HSP_D_R_Q_R 0.1
`define LD5HSP_D_G_HOLD_posedge_negedge 0.1
`define LD5HSP_D_G_HOLD_negedge_negedge 0.1
`define LD5HSP_D_G_SETUP_posedge_negedge 0.1
`define LD5HSP_D_G_SETUP_negedge_negedge 0.1
`define LD5HSP_G_PWH 0.1
`define LD5HSP_SD_PWL 0.1
`define LD5HSP_SD_G_REC_posedge_negedge 0.1
`define LD5HSP_SD_G_REM_posedge_negedge 0.1

module LD5HSP (Q, QN, D, G, SD);

   output Q;
   output QN;
   input D;
   input G;
   input SD;


   reg Notifier;


   U_LD_P_SN_NOTI u0 (IQ, D, G, SD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   not  (GX, G);
   not  (D_, D);
   specify
`ifdef verifault

      if (G && SD) (D -=> QN) = (`LD5HSP_D_F_QN_R,`LD5HSP_D_R_QN_F);
      if (G && SD) (D +=> Q) = (`LD5HSP_D_R_Q_R,`LD5HSP_D_F_Q_F);
      if(SD) (posedge G => (Q +: D)) = (`LD5HSP_G_R_Q_R, `LD5HSP_G_R_Q_F);
      if(SD) (posedge G => (QN -: D)) = (`LD5HSP_G_R_QN_R, `LD5HSP_G_R_QN_F);
      if(!D && G) (posedge SD => (Q +: 1'b0)) = (`LD5HSP_SD_F_Q_R,`LD5HSP_SD_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`LD5HSP_SD_F_Q_R,`LD5HSP_SD_R_Q_F);
      if(!D && G) (posedge SD => (QN +: 1'b1)) = (`LD5HSP_SD_R_QN_R,`LD5HSP_SD_F_QN_F);
      (negedge SD => (QN +: 1'b0)) = (`LD5HSP_SD_R_QN_R,`LD5HSP_SD_F_QN_F);

	$setuphold(negedge G &&& SD, posedge D, `LD5HSP_D_G_SETUP_posedge_negedge, `LD5HSP_D_G_HOLD_posedge_negedge, Notifier);
	$setuphold(negedge G &&& SD, negedge D, `LD5HSP_D_G_SETUP_negedge_negedge, `LD5HSP_D_G_HOLD_negedge_negedge, Notifier);

      $width(posedge G, `LD5HSP_G_PWH, 0, Notifier);
      $width(negedge SD, `LD5HSP_SD_PWL, 0, Notifier);
	$recovery(posedge SD, negedge G &&& D_, `LD5HSP_SD_G_REC_posedge_negedge, Notifier);

	$hold(negedge G &&& D_, posedge SD, `LD5HSP_SD_G_REM_posedge_negedge, Notifier);
`else

      (D -=> QN) = (`LD5HSP_D_F_QN_R,`LD5HSP_D_R_QN_F);
      (D +=> Q) = (`LD5HSP_D_R_Q_R,`LD5HSP_D_F_Q_F);
      (posedge G => (Q +: D)) = (`LD5HSP_G_R_Q_R, `LD5HSP_G_R_Q_F);
            (posedge G => (QN -: D)) = (`LD5HSP_G_R_QN_R, `LD5HSP_G_R_QN_F);
      (posedge SD => (Q +: 1'b0)) = (`LD5HSP_SD_F_Q_R,`LD5HSP_SD_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`LD5HSP_SD_F_Q_R,`LD5HSP_SD_R_Q_F);
      (posedge SD => (QN +: 1'b1)) = (`LD5HSP_SD_R_QN_R,`LD5HSP_SD_F_QN_F);
      (negedge SD => (QN +: 1'b0)) = (`LD5HSP_SD_R_QN_R,`LD5HSP_SD_F_QN_F);
 
        $setuphold(negedge G &&& SD, posedge D, `LD5HSP_D_G_SETUP_posedge_negedge, `LD5HSP_D_G_HOLD_posedge_negedge, Notifier);
        $setuphold(negedge G &&& SD, negedge D, `LD5HSP_D_G_SETUP_negedge_negedge, `LD5HSP_D_G_HOLD_negedge_negedge, Notifier);
 
      $width(posedge G, `LD5HSP_G_PWH, 0, Notifier);
      $width(negedge SD, `LD5HSP_SD_PWL, 0, Notifier);
        $recovery(posedge SD, negedge G &&& D_, `LD5HSP_SD_G_REC_posedge_negedge, Notifier);
 
        $hold(negedge G &&& D_, posedge SD, `LD5HSP_SD_G_REM_posedge_negedge, Notifier);

`endif
   endspecify
`endif


endmodule // LD5HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:27 and Version :1.1 //
 
//  START 
// CELL LD6HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD6HS_SD_F_QN_F 0.1
`define LD6HS_SD_R_QN_R 0.1
`define LD6HS_GN_F_QN_F 0.1
`define LD6HS_GN_F_QN_R 0.1
`define LD6HS_D_F_QN_R 0.1
`define LD6HS_D_R_QN_F 0.1
`define LD6HS_SD_F_Q_R 0.1
`define LD6HS_SD_R_Q_F 0.1
`define LD6HS_GN_F_Q_R 0.1
`define LD6HS_GN_F_Q_F 0.1
`define LD6HS_D_F_Q_F 0.1
`define LD6HS_D_R_Q_R 0.1
`define LD6HS_D_GN_HOLD_posedge_posedge 0.1
`define LD6HS_D_GN_HOLD_negedge_posedge 0.1
`define LD6HS_D_GN_SETUP_posedge_posedge 0.1
`define LD6HS_D_GN_SETUP_negedge_posedge 0.1
`define LD6HS_GN_PWL 0.1
`define LD6HS_SD_PWL 0.1
`define LD6HS_SD_GN_REC_posedge_posedge 0.1
`define LD6HS_SD_GN_REM_posedge_posedge 0.1

module LD6HS (Q, QN, D, GN, SD);

   output Q;
   output QN;
   input D;
   input GN;
   input SD;


   reg Notifier;


   U_LD_N_SN_NOTI u0 (IQ, D, GN, SD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
    not  (D_, D);
 
   specify
`ifdef verifault

      if (!GN && SD) (D -=> QN) = (`LD6HS_D_F_QN_R,`LD6HS_D_R_QN_F);
      if (!GN && SD) (D +=> Q) = (`LD6HS_D_R_Q_R,`LD6HS_D_F_Q_F);
      if(SD) (negedge GN => (Q +: D)) = (`LD6HS_GN_F_Q_R, `LD6HS_GN_F_Q_F);
      if(SD) (negedge GN => (QN -: D)) = (`LD6HS_GN_F_QN_R, `LD6HS_GN_F_QN_F);
      if(!D && !GN) (posedge SD => (Q +: 1'b0)) = (`LD6HS_SD_F_Q_R,`LD6HS_SD_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`LD6HS_SD_F_Q_R,`LD6HS_SD_R_Q_F);
      if(!D && !GN) (posedge SD => (QN +: 1'b1)) = (`LD6HS_SD_R_QN_R,`LD6HS_SD_F_QN_F);
      (negedge SD => (QN +: 1'b0)) = (`LD6HS_SD_R_QN_R,`LD6HS_SD_F_QN_F);

	$setuphold(posedge GN &&& SD, posedge D, `LD6HS_D_GN_SETUP_posedge_posedge, `LD6HS_D_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& SD, negedge D, `LD6HS_D_GN_SETUP_negedge_posedge, `LD6HS_D_GN_HOLD_negedge_posedge, Notifier);

      $width(negedge GN, `LD6HS_GN_PWL, 0, Notifier);
      $width(negedge SD, `LD6HS_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge GN &&& D_, `LD6HS_SD_GN_REC_posedge_posedge, Notifier);

	$hold(posedge GN &&& D_, posedge SD, `LD6HS_SD_GN_REM_posedge_posedge, Notifier);

`else

      (D -=> QN) = (`LD6HS_D_F_QN_R,`LD6HS_D_R_QN_F);
      (D +=> Q) = (`LD6HS_D_R_Q_R,`LD6HS_D_F_Q_F);
      (negedge GN => (Q +: D)) = (`LD6HS_GN_F_Q_R, `LD6HS_GN_F_Q_F);
      (negedge GN => (QN -: D)) = (`LD6HS_GN_F_QN_R, `LD6HS_GN_F_QN_F);
      (posedge SD => (Q +: 1'b0)) = (`LD6HS_SD_F_Q_R,`LD6HS_SD_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`LD6HS_SD_F_Q_R,`LD6HS_SD_R_Q_F);
      (posedge SD => (QN +: 1'b1)) = (`LD6HS_SD_R_QN_R,`LD6HS_SD_F_QN_F);
      (negedge SD => (QN +: 1'b0)) = (`LD6HS_SD_R_QN_R,`LD6HS_SD_F_QN_F);
 
        $setuphold(posedge GN &&& SD, posedge D, `LD6HS_D_GN_SETUP_posedge_posedge, `LD6HS_D_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& SD, negedge D, `LD6HS_D_GN_SETUP_negedge_posedge, `LD6HS_D_GN_HOLD_negedge_posedge, Notifier);
 
      $width(negedge GN, `LD6HS_GN_PWL, 0, Notifier);
      $width(negedge SD, `LD6HS_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge GN &&& D_, `LD6HS_SD_GN_REC_posedge_posedge, Notifier);
 
        $hold(posedge GN &&& D_, posedge SD, `LD6HS_SD_GN_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD6HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:30 and Version :1.1 //
 
//  START 
// CELL LD6HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD6HSP_SD_F_QN_F 0.1
`define LD6HSP_SD_R_QN_R 0.1
`define LD6HSP_GN_F_QN_F 0.1
`define LD6HSP_GN_F_QN_R 0.1
`define LD6HSP_D_F_QN_R 0.1
`define LD6HSP_D_R_QN_F 0.1
`define LD6HSP_SD_F_Q_R 0.1
`define LD6HSP_SD_R_Q_F 0.1
`define LD6HSP_GN_F_Q_R 0.1
`define LD6HSP_GN_F_Q_F 0.1
`define LD6HSP_D_F_Q_F 0.1
`define LD6HSP_D_R_Q_R 0.1
`define LD6HSP_D_GN_HOLD_posedge_posedge 0.1
`define LD6HSP_D_GN_HOLD_negedge_posedge 0.1
`define LD6HSP_D_GN_SETUP_posedge_posedge 0.1
`define LD6HSP_D_GN_SETUP_negedge_posedge 0.1
`define LD6HSP_GN_PWL 0.1
`define LD6HSP_SD_PWL 0.1
`define LD6HSP_SD_GN_REC_posedge_posedge 0.1
`define LD6HSP_SD_GN_REM_posedge_posedge 0.1

module LD6HSP (Q, QN, D, GN, SD);

   output Q;
   output QN;
   input D;
   input GN;
   input SD;


   reg Notifier;


   U_LD_N_SN_NOTI u0 (IQ, D, GN, SD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
    not  (D_, D);
 
   specify
`ifdef verifault

      if (!GN && SD) (D -=> QN) = (`LD6HSP_D_F_QN_R,`LD6HSP_D_R_QN_F);
      if (!GN && SD) (D +=> Q) = (`LD6HSP_D_R_Q_R,`LD6HSP_D_F_Q_F);
      if(SD) (negedge GN => (Q +: D)) = (`LD6HSP_GN_F_Q_R, `LD6HSP_GN_F_Q_F);
      if(SD) (negedge GN => (QN -: D)) = (`LD6HSP_GN_F_QN_R, `LD6HSP_GN_F_QN_F);
      if(!D && !GN) (posedge SD => (Q +: 1'b0)) = (`LD6HSP_SD_F_Q_R,`LD6HSP_SD_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`LD6HSP_SD_F_Q_R,`LD6HSP_SD_R_Q_F);
      if(!D && !GN) (posedge SD => (QN +: 1'b1)) = (`LD6HSP_SD_R_QN_R,`LD6HSP_SD_F_QN_F);
      (negedge SD => (QN +: 1'b0)) = (`LD6HSP_SD_R_QN_R,`LD6HSP_SD_F_QN_F);

	$setuphold(posedge GN &&& SD, posedge D, `LD6HSP_D_GN_SETUP_posedge_posedge, `LD6HSP_D_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& SD, negedge D, `LD6HSP_D_GN_SETUP_negedge_posedge, `LD6HSP_D_GN_HOLD_negedge_posedge, Notifier);

      $width(negedge GN, `LD6HSP_GN_PWL, 0, Notifier);
      $width(negedge SD, `LD6HSP_SD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge GN &&& D_, `LD6HSP_SD_GN_REC_posedge_posedge, Notifier);

	$hold(posedge GN &&& D_, posedge SD, `LD6HSP_SD_GN_REM_posedge_posedge, Notifier);

`else

      (D -=> QN) = (`LD6HSP_D_F_QN_R,`LD6HSP_D_R_QN_F);
      (D +=> Q) = (`LD6HSP_D_R_Q_R,`LD6HSP_D_F_Q_F);
      (negedge GN => (Q +: D)) = (`LD6HSP_GN_F_Q_R, `LD6HSP_GN_F_Q_F);
      (negedge GN => (QN -: D)) = (`LD6HSP_GN_F_QN_R, `LD6HSP_GN_F_QN_F);
      (posedge SD => (Q +: 1'b0)) = (`LD6HSP_SD_F_Q_R,`LD6HSP_SD_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`LD6HSP_SD_F_Q_R,`LD6HSP_SD_R_Q_F);
      (posedge SD => (QN +: 1'b1)) = (`LD6HSP_SD_R_QN_R,`LD6HSP_SD_F_QN_F);
      (negedge SD => (QN +: 1'b0)) = (`LD6HSP_SD_R_QN_R,`LD6HSP_SD_F_QN_F);
 
        $setuphold(posedge GN &&& SD, posedge D, `LD6HSP_D_GN_SETUP_posedge_posedge, `LD6HSP_D_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& SD, negedge D, `LD6HSP_D_GN_SETUP_negedge_posedge, `LD6HSP_D_GN_HOLD_negedge_posedge, Notifier);
 
      $width(negedge GN, `LD6HSP_GN_PWL, 0, Notifier);
      $width(negedge SD, `LD6HSP_SD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge GN &&& D_, `LD6HSP_SD_GN_REC_posedge_posedge, Notifier);
 
        $hold(posedge GN &&& D_, posedge SD, `LD6HSP_SD_GN_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD6HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:30 and Version :1.1 //
 
//  START 
// CELL LD7HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD7HS_SD_F_QN_F 0.1
`define LD7HS_SD_R_QN_R 0.1
`define LD7HS_CD_F_QN_R 0.1
`define LD7HS_CD_R_QN_F 0.1
`define LD7HS_GN_F_QN_F 0.1
`define LD7HS_GN_F_QN_R 0.1
`define LD7HS_D_F_QN_R 0.1
`define LD7HS_D_R_QN_F 0.1
`define LD7HS_SD_F_Q_R 0.1
`define LD7HS_SD_R_Q_F 0.1
`define LD7HS_CD_F_Q_F 0.1
`define LD7HS_CD_R_Q_R 0.1
`define LD7HS_GN_F_Q_R 0.1
`define LD7HS_GN_F_Q_F 0.1
`define LD7HS_D_F_Q_F 0.1
`define LD7HS_D_R_Q_R 0.1
`define LD7HS_D_GN_HOLD_posedge_posedge 0.1
`define LD7HS_D_GN_HOLD_negedge_posedge 0.1
`define LD7HS_D_GN_SETUP_posedge_posedge 0.1
`define LD7HS_D_GN_SETUP_negedge_posedge 0.1
`define LD7HS_GN_PWL 0.1
`define LD7HS_SD_PWL 0.1
`define LD7HS_CD_PWL 0.1
`define LD7HS_SD_GN_REC_posedge_posedge 0.1
`define LD7HS_CD_GN_REC_posedge_posedge 0.1
`define LD7HS_SD_GN_REM_posedge_posedge 0.1
`define LD7HS_CD_GN_REM_posedge_posedge 0.1
`define LD7HS_SD_CD_REC_posedge_posedge 0.1
`define LD7HS_SD_CD_REM_posedge_posedge 0.1

module LD7HS (Q, QN, D, GN, CD, SD);

   output Q;
   output QN;
   input D;
   input GN;
   input CD;
   input SD;


   reg Notifier;


   U_LD_N_RN_SN_NOTI u0 (IQ, D, GN, CD, SD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   and  (AndGNSD_, GN, SD);
   and  (AndGNCD_, GN, CD);
   and  (AndCDSD_, CD, SD);
   and  (AndSDD, SD, D);
   not  (D_, D);
   and  (AndCDD_, CD, D_);

   specify
`ifdef verifault

      if (!GN && CD && SD) (D -=> QN) = (`LD7HS_D_F_QN_R,`LD7HS_D_R_QN_F);
      if (!GN && CD && SD) (D +=> Q) = (`LD7HS_D_R_Q_R,`LD7HS_D_F_Q_F);
      if(SD && CD) (negedge GN => (Q +: D)) = (`LD7HS_GN_F_Q_R, `LD7HS_GN_F_Q_F);
      if(SD && CD) (negedge GN => (QN -: D)) = (`LD7HS_GN_F_QN_R, `LD7HS_GN_F_QN_F);
      if(D && !GN && SD) (posedge CD => (Q +: 1'b1)) = (`LD7HS_CD_R_Q_R,`LD7HS_CD_F_Q_F);
      if(D && SD || GN && SD) (negedge CD => (Q +: 1'b0)) = (`LD7HS_CD_R_Q_R,`LD7HS_CD_F_Q_F);
      if(!CD || !D && !GN) (posedge SD => (Q +: 1'b0)) = (`LD7HS_SD_F_Q_R,`LD7HS_SD_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`LD7HS_SD_F_Q_R,`LD7HS_SD_R_Q_F);
      if(D && !GN && SD) (posedge CD => (QN +: 1'b0)) = (`LD7HS_CD_F_QN_R,`LD7HS_CD_R_QN_F);
      if(D && SD || GN && SD) (negedge CD => (QN +: 1'b1)) = (`LD7HS_CD_F_QN_R,`LD7HS_CD_R_QN_F);
      if(!CD || !D && !GN) (posedge SD => (QN +: 1'b1)) = (`LD7HS_SD_R_QN_R,`LD7HS_SD_F_QN_F);
      (negedge SD => (QN +: 1'b0)) = (`LD7HS_SD_R_QN_R,`LD7HS_SD_F_QN_F);

	$setuphold(posedge GN &&& AndCDSD_, posedge D, `LD7HS_D_GN_SETUP_posedge_posedge, `LD7HS_D_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& AndCDSD_, negedge D, `LD7HS_D_GN_SETUP_negedge_posedge, `LD7HS_D_GN_HOLD_negedge_posedge, Notifier);

      $width(negedge GN, `LD7HS_GN_PWL, 0, Notifier);
      $width(negedge SD, `LD7HS_SD_PWL, 0, Notifier);
      $width(negedge CD, `LD7HS_CD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge GN &&& AndCDD_, `LD7HS_SD_GN_REC_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge GN &&& AndSDD, `LD7HS_CD_GN_REC_posedge_posedge, Notifier);

	$hold(posedge GN &&& AndCDD_, posedge SD, `LD7HS_SD_GN_REM_posedge_posedge, Notifier);

	$hold(posedge GN &&& AndSDD, posedge CD, `LD7HS_CD_GN_REM_posedge_posedge, Notifier);

	$recovery(posedge SD, posedge CD, `LD7HS_SD_CD_REC_posedge_posedge, Notifier);

	$hold(posedge CD, posedge SD, `LD7HS_SD_CD_REM_posedge_posedge, Notifier);

`else


      (D -=> QN) = (`LD7HS_D_F_QN_R,`LD7HS_D_R_QN_F);
      (D +=> Q) = (`LD7HS_D_R_Q_R,`LD7HS_D_F_Q_F);
      (negedge GN => (Q +: D)) = (`LD7HS_GN_F_Q_R, `LD7HS_GN_F_Q_F);
      (negedge GN => (QN -: D)) = (`LD7HS_GN_F_QN_R, `LD7HS_GN_F_QN_F);
      (posedge CD => (Q +: 1'b1)) = (`LD7HS_CD_R_Q_R,`LD7HS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD7HS_CD_R_Q_R,`LD7HS_CD_F_Q_F);
      (posedge SD => (Q +: 1'b0)) = (`LD7HS_SD_F_Q_R,`LD7HS_SD_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`LD7HS_SD_F_Q_R,`LD7HS_SD_R_Q_F);
      (posedge CD => (QN +: 1'b0)) = (`LD7HS_CD_F_QN_R,`LD7HS_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`LD7HS_CD_F_QN_R,`LD7HS_CD_R_QN_F);
      (posedge SD => (QN +: 1'b1)) = (`LD7HS_SD_R_QN_R,`LD7HS_SD_F_QN_F);
      (negedge SD => (QN +: 1'b0)) = (`LD7HS_SD_R_QN_R,`LD7HS_SD_F_QN_F);
 
        $setuphold(posedge GN &&& AndCDSD_, posedge D, `LD7HS_D_GN_SETUP_posedge_posedge, `LD7HS_D_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& AndCDSD_, negedge D, `LD7HS_D_GN_SETUP_negedge_posedge, `LD7HS_D_GN_HOLD_negedge_posedge, Notifier);
 
      $width(negedge GN, `LD7HS_GN_PWL, 0, Notifier);
      $width(negedge SD, `LD7HS_SD_PWL, 0, Notifier);
      $width(negedge CD, `LD7HS_CD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge GN &&& AndCDD_, `LD7HS_SD_GN_REC_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge GN &&& AndSDD, `LD7HS_CD_GN_REC_posedge_posedge, Notifier);
 
        $hold(posedge GN &&& AndCDD_, posedge SD, `LD7HS_SD_GN_REM_posedge_posedge, Notifier);
 
        $hold(posedge GN &&& AndSDD, posedge CD, `LD7HS_CD_GN_REM_posedge_posedge, Notifier);
 
        $recovery(posedge SD, posedge CD, `LD7HS_SD_CD_REC_posedge_posedge, Notifier);
 
        $hold(posedge CD, posedge SD, `LD7HS_SD_CD_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD7HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:34 and Version :1.1 //
 
//  START 
// CELL LD7HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LD7HSP_SD_F_QN_F 0.1
`define LD7HSP_SD_R_QN_R 0.1
`define LD7HSP_CD_F_QN_R 0.1
`define LD7HSP_CD_R_QN_F 0.1
`define LD7HSP_GN_F_QN_F 0.1
`define LD7HSP_GN_F_QN_R 0.1
`define LD7HSP_D_F_QN_R 0.1
`define LD7HSP_D_R_QN_F 0.1
`define LD7HSP_SD_F_Q_R 0.1
`define LD7HSP_SD_R_Q_F 0.1
`define LD7HSP_CD_F_Q_F 0.1
`define LD7HSP_CD_R_Q_R 0.1
`define LD7HSP_GN_F_Q_R 0.1
`define LD7HSP_GN_F_Q_F 0.1
`define LD7HSP_D_F_Q_F 0.1
`define LD7HSP_D_R_Q_R 0.1
`define LD7HSP_D_GN_HOLD_posedge_posedge 0.1
`define LD7HSP_D_GN_HOLD_negedge_posedge 0.1
`define LD7HSP_D_GN_SETUP_posedge_posedge 0.1
`define LD7HSP_D_GN_SETUP_negedge_posedge 0.1
`define LD7HSP_GN_PWL 0.1
`define LD7HSP_SD_PWL 0.1
`define LD7HSP_CD_PWL 0.1
`define LD7HSP_SD_GN_REC_posedge_posedge 0.1
`define LD7HSP_CD_GN_REC_posedge_posedge 0.1
`define LD7HSP_SD_GN_REM_posedge_posedge 0.1
`define LD7HSP_CD_GN_REM_posedge_posedge 0.1
`define LD7HSP_SD_CD_REC_posedge_posedge 0.1
`define LD7HSP_SD_CD_REM_posedge_posedge 0.1

module LD7HSP (Q, QN, D, GN, CD, SD);

   output Q;
   output QN;
   input D;
   input GN;
   input CD;
   input SD;


   reg Notifier;


   U_LD_N_RN_SN_NOTI u0 (IQ, D, GN, CD, SD, Notifier);

   buf  u1 (Q, IQ);
   not  u2 (QN, IQ);



`ifdef functional
`else
   and  (AndGNSD_, GN, SD);
   and  (AndGNCD_, GN, CD);
   and  (AndCDSD_, CD, SD);
   and  (AndSDD, SD, D);
   not  (D_, D);
   and  (AndCDD_, CD, D_);

   specify
`ifdef verifault

      if (!GN && CD && SD) (D -=> QN) = (`LD7HSP_D_F_QN_R,`LD7HSP_D_R_QN_F);
      if (!GN && CD && SD) (D +=> Q) = (`LD7HSP_D_R_Q_R,`LD7HSP_D_F_Q_F);
      if(SD && CD) (negedge GN => (Q +: D)) = (`LD7HSP_GN_F_Q_R, `LD7HSP_GN_F_Q_F);
      if(SD && CD) (negedge GN => (QN -: D)) = (`LD7HSP_GN_F_QN_R, `LD7HSP_GN_F_QN_F);
      if(D && !GN && SD) (posedge CD => (Q +: 1'b1)) = (`LD7HSP_CD_R_Q_R,`LD7HSP_CD_F_Q_F);
      if(D && SD || GN && SD) (negedge CD => (Q +: 1'b0)) = (`LD7HSP_CD_R_Q_R,`LD7HSP_CD_F_Q_F);
      if(!CD || !D && !GN) (posedge SD => (Q +: 1'b0)) = (`LD7HSP_SD_F_Q_R,`LD7HSP_SD_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`LD7HSP_SD_F_Q_R,`LD7HSP_SD_R_Q_F);
      if(D && !GN && SD) (posedge CD => (QN +: 1'b0)) = (`LD7HSP_CD_F_QN_R,`LD7HSP_CD_R_QN_F);
      if(D && SD || GN && SD) (negedge CD => (QN +: 1'b1)) = (`LD7HSP_CD_F_QN_R,`LD7HSP_CD_R_QN_F);
      if(!CD || !D && !GN) (posedge SD => (QN +: 1'b1)) = (`LD7HSP_SD_R_QN_R,`LD7HSP_SD_F_QN_F);
      (negedge SD => (QN +: 1'b0)) = (`LD7HSP_SD_R_QN_R,`LD7HSP_SD_F_QN_F);

	$setuphold(posedge GN &&& AndCDSD_, posedge D, `LD7HSP_D_GN_SETUP_posedge_posedge, `LD7HSP_D_GN_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge GN &&& AndCDSD_, negedge D, `LD7HSP_D_GN_SETUP_negedge_posedge, `LD7HSP_D_GN_HOLD_negedge_posedge, Notifier);

      $width(negedge GN, `LD7HSP_GN_PWL, 0, Notifier);
      $width(negedge SD, `LD7HSP_SD_PWL, 0, Notifier);
      $width(negedge CD, `LD7HSP_CD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge GN &&& AndCDD_, `LD7HSP_SD_GN_REC_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge GN &&& AndSDD, `LD7HSP_CD_GN_REC_posedge_posedge, Notifier);

	$hold(posedge GN &&& AndCDD_, posedge SD, `LD7HSP_SD_GN_REM_posedge_posedge, Notifier);

	$hold(posedge GN &&& AndSDD, posedge CD, `LD7HSP_CD_GN_REM_posedge_posedge, Notifier);

	$recovery(posedge SD, posedge CD, `LD7HSP_SD_CD_REC_posedge_posedge, Notifier);

	$hold(posedge CD, posedge SD, `LD7HSP_SD_CD_REM_posedge_posedge, Notifier);

`else


      (D -=> QN) = (`LD7HSP_D_F_QN_R,`LD7HSP_D_R_QN_F);
      (D +=> Q) = (`LD7HSP_D_R_Q_R,`LD7HSP_D_F_Q_F);
      (negedge GN => (Q +: D)) = (`LD7HSP_GN_F_Q_R, `LD7HSP_GN_F_Q_F);
      (negedge GN => (QN -: D)) = (`LD7HSP_GN_F_QN_R, `LD7HSP_GN_F_QN_F);
      (posedge CD => (Q +: 1'b1)) = (`LD7HSP_CD_R_Q_R,`LD7HSP_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`LD7HSP_CD_R_Q_R,`LD7HSP_CD_F_Q_F);
      (posedge SD => (Q +: 1'b0)) = (`LD7HSP_SD_F_Q_R,`LD7HSP_SD_R_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`LD7HSP_SD_F_Q_R,`LD7HSP_SD_R_Q_F);
      (posedge CD => (QN +: 1'b0)) = (`LD7HSP_CD_F_QN_R,`LD7HSP_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`LD7HSP_CD_F_QN_R,`LD7HSP_CD_R_QN_F);
      (posedge SD => (QN +: 1'b1)) = (`LD7HSP_SD_R_QN_R,`LD7HSP_SD_F_QN_F);
      (negedge SD => (QN +: 1'b0)) = (`LD7HSP_SD_R_QN_R,`LD7HSP_SD_F_QN_F);
 
        $setuphold(posedge GN &&& AndCDSD_, posedge D, `LD7HSP_D_GN_SETUP_posedge_posedge, `LD7HSP_D_GN_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge GN &&& AndCDSD_, negedge D, `LD7HSP_D_GN_SETUP_negedge_posedge, `LD7HSP_D_GN_HOLD_negedge_posedge, Notifier);
 
      $width(negedge GN, `LD7HSP_GN_PWL, 0, Notifier);
      $width(negedge SD, `LD7HSP_SD_PWL, 0, Notifier);
      $width(negedge CD, `LD7HSP_CD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge GN &&& AndCDD_, `LD7HSP_SD_GN_REC_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge GN &&& AndSDD, `LD7HSP_CD_GN_REC_posedge_posedge, Notifier);
 
        $hold(posedge GN &&& AndCDD_, posedge SD, `LD7HSP_SD_GN_REM_posedge_posedge, Notifier);
 
        $hold(posedge GN &&& AndSDD, posedge CD, `LD7HSP_CD_GN_REM_posedge_posedge, Notifier);
 
        $recovery(posedge SD, posedge CD, `LD7HSP_SD_CD_REC_posedge_posedge, Notifier);
 
        $hold(posedge CD, posedge SD, `LD7HSP_SD_CD_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule // LD7HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:34 and Version :1.1 //
 
//  START 
// CELL LR1QHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define LR1QHS_SN_F_Q_R 0.1
`define LR1QHS_RN_F_Q_F 0.1
`define LR1QHS_RN_R_Q_R 0.1
`define LR1QHS_RN_SN_REM_posedge_posedge 0.1
`define LR1QHS_RN_SN_REC_posedge_posedge 0.1
`define LR1QHS_RN_PWL 0.1
`define LR1QHS_SN_PWL 0.1

module LR1QHS (Q, RN, SN);

   output Q;
   input RN;
   input SN;


   reg Notifier;


   U_RS_RN_SN_NOTI u0 (   // Verilog Seq UDP
      IQ, RN, SN, Notifier);

   buf  u1 (Q, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      if(!SN)(posedge RN => (Q +: 1'b1)) = (`LR1QHS_RN_R_Q_R,`LR1QHS_RN_F_Q_F);
      (negedge RN => (Q +: 1'b0)) = (`LR1QHS_RN_R_Q_R,`LR1QHS_RN_F_Q_F);
     if(RN) (negedge SN => (Q +: 1'b1)) = (`LR1QHS_SN_F_Q_R,`LR1QHS_SN_F_Q_R);

      $width(negedge SN, `LR1QHS_SN_PWL, 0, Notifier);
      $width(negedge RN, `LR1QHS_RN_PWL, 0, Notifier);
	$recovery(posedge RN, posedge SN, `LR1QHS_RN_SN_REC_posedge_posedge, Notifier);

	$hold(posedge SN, posedge RN, `LR1QHS_RN_SN_REM_posedge_posedge, Notifier);

`else

       (posedge RN => (Q +: 1'b1)) = (`LR1QHS_RN_R_Q_R,`LR1QHS_RN_F_Q_F);
      (negedge RN => (Q +: 1'b0)) = (`LR1QHS_RN_R_Q_R,`LR1QHS_RN_F_Q_F);
       (negedge SN => (Q +: 1'b1)) = (`LR1QHS_SN_F_Q_R,`LR1QHS_SN_F_Q_R);
 
      $width(negedge SN, `LR1QHS_SN_PWL, 0, Notifier);
      $width(negedge RN, `LR1QHS_RN_PWL, 0, Notifier);
        $recovery(posedge RN, posedge SN, `LR1QHS_RN_SN_REC_posedge_posedge, Notifier);
 
        $hold(posedge SN, posedge RN, `LR1QHS_RN_SN_REM_posedge_posedge, Notifier);
`endif
   endspecify
`endif


endmodule
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:47 and Version :1.1 //
 
//  START
 
// CELL MUX21HSX05 

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define MUX21HSX05_S_F_Z_F 0.1
`define MUX21HSX05_S_R_Z_R 0.1
`define MUX21HSX05_S_F_Z_R 0.1
`define MUX21HSX05_S_R_Z_F 0.1
`define MUX21HSX05_B_F_Z_F 0.1
`define MUX21HSX05_B_R_Z_R 0.1
`define MUX21HSX05_A_F_Z_F 0.1
`define MUX21HSX05_A_R_Z_R 0.1

module MUX21HSX05 (Z, A, B, S);

   output Z;
   input A;
   input B;
   input S;


   U_MUX2  u0 (Z, A, B, S);

   buf u1 (ST, S);
   buf u2 (BT, B);
   buf u3 (AT, A);
 
`ifdef tristatecheck
always @(ST or AT or BT)
  begin
        if (((B === 1'bz) && (S == 1)) || ((A === 1'bz) && (S == 0)) || ((S === 1'bx) && ((A === 1'bz) || (B === 1'bz))))
        $display ("WARNING: Cell MUX21HSX05 used in IDDQ unsafe mode with A = %b, B = %b, S = %b at time %d", A, B, S,$time);
  end
`endif


`ifdef functional
`else
   specify

      if (!A && B) (S +=> Z) = (`MUX21HSX05_S_R_Z_R,`MUX21HSX05_S_F_Z_F);
      if (A && !B) (S -=> Z) = (`MUX21HSX05_S_F_Z_R,`MUX21HSX05_S_R_Z_F);
      (B +=> Z) = (`MUX21HSX05_B_R_Z_R,`MUX21HSX05_B_F_Z_F);
      (A +=> Z) = (`MUX21HSX05_A_R_Z_R,`MUX21HSX05_A_F_Z_F);

   endspecify
`endif


endmodule // MUX21HSX05

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
//  END
// Created from CVS on Date :1998/07/07 13:18:59 and Version :1.1 //
 
//  START
// CELL MUX21HS 

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define MUX21HS_S_F_Z_F 0.1
`define MUX21HS_S_R_Z_R 0.1
`define MUX21HS_S_F_Z_R 0.1
`define MUX21HS_S_R_Z_F 0.1
`define MUX21HS_B_F_Z_F 0.1
`define MUX21HS_B_R_Z_R 0.1
`define MUX21HS_A_F_Z_F 0.1
`define MUX21HS_A_R_Z_R 0.1

module MUX21HS (Z, A, B, S);

   output Z;
   input A;
   input B;
   input S;


   U_MUX2  u0 (Z, A, B, S);

   buf u1 (ST, S);
   buf u2 (BT, B);
   buf u3 (AT, A);
 
`ifdef tristatecheck
always @(ST or AT or BT)
  begin
        if (((B === 1'bz) && (S == 1)) || ((A === 1'bz) && (S == 0)) || ((S === 1'bx) && ((A === 1'bz) || (B === 1'bz))))
        $display ("WARNING: Cell MUX21HS used in IDDQ unsafe mode with A = %b, B = %b, S = %b at time %d", A, B, S,$time);
  end
`endif


`ifdef functional
`else
   specify

      if (!A && B) (S +=> Z) = (`MUX21HS_S_R_Z_R,`MUX21HS_S_F_Z_F);
      if (A && !B) (S -=> Z) = (`MUX21HS_S_F_Z_R,`MUX21HS_S_R_Z_F);
      (B +=> Z) = (`MUX21HS_B_R_Z_R,`MUX21HS_B_F_Z_F);
      (A +=> Z) = (`MUX21HS_A_R_Z_R,`MUX21HS_A_F_Z_F);

   endspecify
`endif


endmodule // MUX21HS

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
//  END
// Created from CVS on Date :1998/07/07 13:18:59 and Version :1.1 //
 
//  START
// CELL MUX21HSP 

`celldefine
`define functional //off sdf
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define MUX21HSP_S_F_Z_F 0.1
`define MUX21HSP_S_R_Z_R 0.1
`define MUX21HSP_S_F_Z_R 0.1
`define MUX21HSP_S_R_Z_F 0.1
`define MUX21HSP_B_F_Z_F 0.1
`define MUX21HSP_B_R_Z_R 0.1
`define MUX21HSP_A_F_Z_F 0.1
`define MUX21HSP_A_R_Z_R 0.1

module MUX21HSP (Z, A, B, S);

   output Z;
   input A;
   input B;
   input S;


   U_MUX2  u0 (Z, A, B, S);

   buf u1 (ST, S);
   buf u2 (BT, B);
   buf u3 (AT, A);
 
`ifdef tristatecheck
always @(ST or AT or BT)
  begin
        if (((B === 1'bz) && (S == 1)) || ((A === 1'bz) && (S == 0)) || ((S === 1'bx) && ((A === 1'bz) || (B === 1'bz))))
        $display ("WARNING: Cell MUX21HSP used in IDDQ unsafe mode with A = %b, B = %b, S = %b at time %d", A, B, S,$time);
  end
`endif


`ifdef functional
`else
   specify

      if (!A && B) (S +=> Z) = (`MUX21HSP_S_R_Z_R,`MUX21HSP_S_F_Z_F);
      if (A && !B) (S -=> Z) = (`MUX21HSP_S_F_Z_R,`MUX21HSP_S_R_Z_F);
      (B +=> Z) = (`MUX21HSP_B_R_Z_R,`MUX21HSP_B_F_Z_F);
      (A +=> Z) = (`MUX21HSP_A_R_Z_R,`MUX21HSP_A_F_Z_F);

   endspecify
`endif


endmodule // MUX21HSP

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
//  END
// Created from CVS on Date :1998/07/07 13:18:59 and Version :1.1 //
 
//  START
// CELL MUX21HSX4 

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define MUX21HSX4_S_F_Z_F 0.1
`define MUX21HSX4_S_R_Z_R 0.1
`define MUX21HSX4_S_F_Z_R 0.1
`define MUX21HSX4_S_R_Z_F 0.1
`define MUX21HSX4_B_F_Z_F 0.1
`define MUX21HSX4_B_R_Z_R 0.1
`define MUX21HSX4_A_F_Z_F 0.1
`define MUX21HSX4_A_R_Z_R 0.1

module MUX21HSX4 (Z, A, B, S);

   output Z;
   input A;
   input B;
   input S;


   U_MUX2  u0 (Z, A, B, S);

   buf u1 (ST, S);
   buf u2 (BT, B);
   buf u3 (AT, A);
 
`ifdef tristatecheck
always @(ST or AT or BT)
  begin
        if (((B === 1'bz) && (S == 1)) || ((A === 1'bz) && (S == 0)) || ((S === 1'bx) && ((A === 1'bz) || (B === 1'bz))))
        $display ("WARNING: Cell MUX21HSX4 used in IDDQ unsafe mode with A = %b, B = %b, S = %b at time %d", A, B, S,$time);
  end
`endif


`ifdef functional
`else
   specify

      if (!A && B) (S +=> Z) = (`MUX21HSX4_S_R_Z_R,`MUX21HSX4_S_F_Z_F);
      if (A && !B) (S -=> Z) = (`MUX21HSX4_S_F_Z_R,`MUX21HSX4_S_R_Z_F);
      (B +=> Z) = (`MUX21HSX4_B_R_Z_R,`MUX21HSX4_B_F_Z_F);
      (A +=> Z) = (`MUX21HSX4_A_R_Z_R,`MUX21HSX4_A_F_Z_F);

   endspecify
`endif


endmodule // MUX21HSX4

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
//  END
// Created from CVS on Date :1998/07/07 13:18:59 and Version :1.1 //
 
//  START
// CELL F_MUX21HSP 

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define F_MUX21HSP_S_F_Z_F 0.1
`define F_MUX21HSP_S_R_Z_R 0.1
`define F_MUX21HSP_S_F_Z_R 0.1
`define F_MUX21HSP_S_R_Z_F 0.1
`define F_MUX21HSP_B_F_Z_F 0.1
`define F_MUX21HSP_B_R_Z_R 0.1
`define F_MUX21HSP_A_F_Z_F 0.1
`define F_MUX21HSP_A_R_Z_R 0.1

module F_MUX21HSP (Z, A, B, S);

   output Z;
   input A;
   input B;
   input S;


   U_MUX2  u0 (Z, A, B, S);

   buf u1 (ST, S);
   buf u2 (BT, B);
   buf u3 (AT, A);
 
`ifdef tristatecheck
always @(ST or AT or BT)
  begin
        if (((B === 1'bz) && (S == 1)) || ((A === 1'bz) && (S == 0)) || ((S === 1'bx) && ((A === 1'bz) || (B === 1'bz))))
        $display ("WARNING: Cell F_MUX21HSP used in IDDQ unsafe mode with A = %b, B = %b, S = %b at time %d", A, B, S,$time);
  end
`endif


`ifdef functional
`else
   specify

      if (!A && B) (S +=> Z) = (`F_MUX21HSP_S_R_Z_R,`F_MUX21HSP_S_F_Z_F);
      if (A && !B) (S -=> Z) = (`F_MUX21HSP_S_F_Z_R,`F_MUX21HSP_S_R_Z_F);
      (B +=> Z) = (`F_MUX21HSP_B_R_Z_R,`F_MUX21HSP_B_F_Z_F);
      (A +=> Z) = (`F_MUX21HSP_A_R_Z_R,`F_MUX21HSP_A_F_Z_F);

   endspecify
`endif


endmodule // F_MUX21HSP

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
//  END
// Created from CVS on Date :1998/07/07 13:18:59 and Version :1.1 //
 
//  START
// Cell MUX21DNHS
 
`celldefine
`ifdef verifault
   `suppress_faults
   `enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 
`define MUX21DNHS_A_R_Z_F 0.1
`define MUX21DNHS_A_F_Z_R 0.1
`define MUX21DNHS_B_R_Z_F 0.1
`define MUX21DNHS_B_F_Z_R 0.1
`define MUX21DNHS_SN_R_Z_R 0.1
`define MUX21DNHS_SN_F_Z_F 0.1
`define MUX21DNHS_SN_R_Z_F 0.1
`define MUX21DNHS_SN_F_Z_R 0.1
`define MUX21DNHS_S_R_Z_R 0.1
`define MUX21DNHS_S_F_Z_F 0.1
`define MUX21DNHS_S_R_Z_F 0.1
`define MUX21DNHS_S_F_Z_R 0.1
 
module MUX21DNHS (Z, A, B, S, SN);
 
        output Z;
        input A;
        input B;
        input S;
        input SN;
 
        tri  ZPREVIOUS;
        not    U1 (INTERNAL4, A) ;
        not    U2 (INTERNAL5, S) ;
        and    U3 (INTERNAL3, INTERNAL4, INTERNAL5) ;
        bufif1    U4 (ZPREVIOUS, 1'b1, INTERNAL3) ;
        nand    U5 (INTERNAL8, A, SN) ;
        bufif0    U6 (ZPREVIOUS, 1'b0, INTERNAL8) ;
        not    U7 (INTERNAL12, B) ;
        not    U8 (INTERNAL13, SN) ;
        and    U9 (INTERNAL11, INTERNAL12, INTERNAL13) ;
        bufif1    U10 (ZPREVIOUS, 1'b1, INTERNAL11) ;
        nand    U11 (INTERNAL16, B, S) ;
        bufif0    U12 (ZPREVIOUS, 1'b0, INTERNAL16) ;
        nmos    U13 (Z, ZPREVIOUS, 1'b1) ;
         
        buf     U14 (ST, S);                                    
        buf     U15 (BT, B);                                    
        buf     U16 (AT, A);                                    
        buf     U17 (SNT,SN); 
`ifdef tristatecheck
always @(ST or SNT or AT or BT)
  begin
        if (((B === 1'bz) && (S == 1) && (SN == 0)) || ((A === 1'bz) && (S == 0) && (SN == 1)) || (((S === 1'bx) || (SN === 1'bx)) && ((A === 1'bz) || (B === 1'bz))))
           $display ("WARNING: Cell MUX21DNHS used in IDDQ unsafe mode with A = %b, B = %b, S = %b, SN = %b at time %d", A , B, S, SN, $time);
  end
`endif
 
`ifdef functional
`else
 
        specify
 
                (A -=> Z) = (`MUX21DNHS_A_F_Z_R,`MUX21DNHS_A_R_Z_F);
                (B -=> Z) = (`MUX21DNHS_B_F_Z_R,`MUX21DNHS_B_R_Z_F);
                if (!A && B) (SN +=> Z) = (`MUX21DNHS_SN_R_Z_R,`MUX21DNHS_SN_F_Z_F);
                if (A && !B) (SN -=> Z) = (`MUX21DNHS_SN_F_Z_R,`MUX21DNHS_SN_R_Z_F);
                if (A && !B) (S +=> Z) = (`MUX21DNHS_S_R_Z_R,`MUX21DNHS_S_F_Z_F);
                if (!A && B) (S -=> Z) = (`MUX21DNHS_S_F_Z_R,`MUX21DNHS_S_R_Z_F);
 
 
        endspecify
 
`endif
 
endmodule // MUX21DNHS
 
`ifdef verifault
   `disable_portfaults
   `nosuppress_faults
`endif
`endcelldefine
// CELL MUX21NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define MUX21NHS_S_F_Z_R 0.1
`define MUX21NHS_S_R_Z_F 0.1
`define MUX21NHS_S_F_Z_F 0.1
`define MUX21NHS_S_R_Z_R 0.1
`define MUX21NHS_B_F_Z_R 0.1
`define MUX21NHS_B_R_Z_F 0.1
`define MUX21NHS_A_F_Z_R 0.1
`define MUX21NHS_A_R_Z_F 0.1

module MUX21NHS (Z, A, B, S);

   output Z;
   input A;
   input B;
   input S;


   not  u0 (AX, A);
   not  u1 (BX, B);
   U_MUX2  u2 (Z, AX, BX, S);


   buf u3 (ST, S);
   buf u4 (BT, B);
   buf u5 (AT, A);
 
`ifdef tristatecheck
always @(ST or AT or BT)
  begin
        if (((B === 1'bz) && (S == 1)) || ((A === 1'bz) && (S == 0)) || ((S === 1'bx) && ((A === 1'bz) || (B === 1'bz))))
        $display ("WARNING: Cell MUX21NHS used in IDDQ unsafe mode with A = %b, B = %b, S = %b at time %d", A, B, S,$time);
  end
`endif

`ifdef functional
`else
   specify

      if (!A && B) (S -=> Z) = (`MUX21NHS_S_F_Z_R,`MUX21NHS_S_R_Z_F);
      if (A && !B) (S +=> Z) = (`MUX21NHS_S_R_Z_R,`MUX21NHS_S_F_Z_F);
      (B -=> Z) = (`MUX21NHS_B_F_Z_R,`MUX21NHS_B_R_Z_F);
      (A -=> Z) = (`MUX21NHS_A_F_Z_R,`MUX21NHS_A_R_Z_F);

   endspecify
`endif


endmodule // MUX21NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:47 and Version :1.1 //
 
//  START 
// CELL MUX21NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define MUX21NHSP_S_F_Z_R 0.1
`define MUX21NHSP_S_R_Z_F 0.1
`define MUX21NHSP_S_F_Z_F 0.1
`define MUX21NHSP_S_R_Z_R 0.1
`define MUX21NHSP_B_F_Z_R 0.1
`define MUX21NHSP_B_R_Z_F 0.1
`define MUX21NHSP_A_F_Z_R 0.1
`define MUX21NHSP_A_R_Z_F 0.1

module MUX21NHSP (Z, A, B, S);

   output Z;
   input A;
   input B;
   input S;


   not  u0 (AX, A);
   not  u1 (BX, B);
   U_MUX2  u2 (Z, AX, BX, S);


   buf u3 (ST, S);
   buf u4 (BT, B);
   buf u5 (AT, A);
 
`ifdef tristatecheck
always @(ST or AT or BT)
  begin
        if (((B === 1'bz) && (S == 1)) || ((A === 1'bz) && (S == 0)) || ((S === 1'bx) && ((A === 1'bz) || (B === 1'bz))))
        $display ("WARNING: Cell MUX21NHSP used in IDDQ unsafe mode with A = %b, B = %b, S = %b at time %d", A, B, S,$time);
  end
`endif

`ifdef functional
`else
   specify

      if (!A && B) (S -=> Z) = (`MUX21NHSP_S_F_Z_R,`MUX21NHSP_S_R_Z_F);
      if (A && !B) (S +=> Z) = (`MUX21NHSP_S_R_Z_R,`MUX21NHSP_S_F_Z_F);
      (B -=> Z) = (`MUX21NHSP_B_F_Z_R,`MUX21NHSP_B_R_Z_F);
      (A -=> Z) = (`MUX21NHSP_A_F_Z_R,`MUX21NHSP_A_R_Z_F);

   endspecify
`endif


endmodule // MUX21NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:47 and Version :1.1 //
 
//  START 
// CELL MUX21NHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define MUX21NHSX4_S_F_Z_R 0.1
`define MUX21NHSX4_S_R_Z_F 0.1
`define MUX21NHSX4_S_F_Z_F 0.1
`define MUX21NHSX4_S_R_Z_R 0.1
`define MUX21NHSX4_B_F_Z_R 0.1
`define MUX21NHSX4_B_R_Z_F 0.1
`define MUX21NHSX4_A_F_Z_R 0.1
`define MUX21NHSX4_A_R_Z_F 0.1

module MUX21NHSX4 (Z, A, B, S);

   output Z;
   input A;
   input B;
   input S;


   not  u0 (AX, A);
   not  u1 (BX, B);
   U_MUX2  u2 (Z, AX, BX, S);


   buf u3 (ST, S);
   buf u4 (BT, B);
   buf u5 (AT, A);
 
`ifdef tristatecheck
always @(ST or AT or BT)
  begin
        if (((B === 1'bz) && (S == 1)) || ((A === 1'bz) && (S == 0)) || ((S === 1'bx) && ((A === 1'bz) || (B === 1'bz))))
        $display ("WARNING: Cell MUX21NHSX4 used in IDDQ unsafe mode with A = %b, B = %b, S = %b at time %d", A, B, S,$time);
  end
`endif

`ifdef functional
`else
   specify

      if (!A && B) (S -=> Z) = (`MUX21NHSX4_S_F_Z_R,`MUX21NHSX4_S_R_Z_F);
      if (A && !B) (S +=> Z) = (`MUX21NHSX4_S_R_Z_R,`MUX21NHSX4_S_F_Z_F);
      (B -=> Z) = (`MUX21NHSX4_B_F_Z_R,`MUX21NHSX4_B_R_Z_F);
      (A -=> Z) = (`MUX21NHSX4_A_F_Z_R,`MUX21NHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // MUX21NHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:47 and Version :1.1 //
 
//  START 
// CELL F_MUX21NHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_MUX21NHS_S_F_Z_R 0.1
`define F_MUX21NHS_S_R_Z_F 0.1
`define F_MUX21NHS_S_F_Z_F 0.1
`define F_MUX21NHS_S_R_Z_R 0.1
`define F_MUX21NHS_B_F_Z_R 0.1
`define F_MUX21NHS_B_R_Z_F 0.1
`define F_MUX21NHS_A_F_Z_R 0.1
`define F_MUX21NHS_A_R_Z_F 0.1

module F_MUX21NHS (Z, A, B, S);

   output Z;
   input A;
   input B;
   input S;


   not  u0 (AX, A);
   not  u1 (BX, B);
   U_MUX2  u2 (Z, AX, BX, S);


   buf u3 (ST, S);
   buf u4 (BT, B);
   buf u5 (AT, A);
 
`ifdef tristatecheck
always @(ST or AT or BT)
  begin
        if (((B === 1'bz) && (S == 1)) || ((A === 1'bz) && (S == 0)) || ((S === 1'bx) && ((A === 1'bz) || (B === 1'bz))))
        $display ("WARNING: Cell F_MUX21NHS used in IDDQ unsafe mode with A = %b, B = %b, S = %b at time %d", A, B, S,$time);
  end
`endif

`ifdef functional
`else
   specify

      if (!A && B) (S -=> Z) = (`F_MUX21NHS_S_F_Z_R,`F_MUX21NHS_S_R_Z_F);
      if (A && !B) (S +=> Z) = (`F_MUX21NHS_S_R_Z_R,`F_MUX21NHS_S_F_Z_F);
      (B -=> Z) = (`F_MUX21NHS_B_F_Z_R,`F_MUX21NHS_B_R_Z_F);
      (A -=> Z) = (`F_MUX21NHS_A_F_Z_R,`F_MUX21NHS_A_R_Z_F);

   endspecify
`endif


endmodule // F_MUX21NHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:47 and Version :1.1 //
 
//  START 
// CELL F_MUX21NHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_MUX21NHSP_S_F_Z_R 0.1
`define F_MUX21NHSP_S_R_Z_F 0.1
`define F_MUX21NHSP_S_F_Z_F 0.1
`define F_MUX21NHSP_S_R_Z_R 0.1
`define F_MUX21NHSP_B_F_Z_R 0.1
`define F_MUX21NHSP_B_R_Z_F 0.1
`define F_MUX21NHSP_A_F_Z_R 0.1
`define F_MUX21NHSP_A_R_Z_F 0.1

module F_MUX21NHSP (Z, A, B, S);

   output Z;
   input A;
   input B;
   input S;


   not  u0 (AX, A);
   not  u1 (BX, B);
   U_MUX2  u2 (Z, AX, BX, S);


   buf u3 (ST, S);
   buf u4 (BT, B);
   buf u5 (AT, A);
 
`ifdef tristatecheck
always @(ST or AT or BT)
  begin
        if (((B === 1'bz) && (S == 1)) || ((A === 1'bz) && (S == 0)) || ((S === 1'bx) && ((A === 1'bz) || (B === 1'bz))))
        $display ("WARNING: Cell F_MUX21NHSP used in IDDQ unsafe mode with A = %b, B = %b, S = %b at time %d", A, B, S,$time);
  end
`endif

`ifdef functional
`else
   specify

      if (!A && B) (S -=> Z) = (`F_MUX21NHSP_S_F_Z_R,`F_MUX21NHSP_S_R_Z_F);
      if (A && !B) (S +=> Z) = (`F_MUX21NHSP_S_R_Z_R,`F_MUX21NHSP_S_F_Z_F);
      (B -=> Z) = (`F_MUX21NHSP_B_F_Z_R,`F_MUX21NHSP_B_R_Z_F);
      (A -=> Z) = (`F_MUX21NHSP_A_F_Z_R,`F_MUX21NHSP_A_R_Z_F);

   endspecify
`endif


endmodule // F_MUX21NHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:47 and Version :1.1 //
 
//  START 
// CELL F_MUX21NHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_MUX21NHSX4_S_F_Z_R 0.1
`define F_MUX21NHSX4_S_R_Z_F 0.1
`define F_MUX21NHSX4_S_F_Z_F 0.1
`define F_MUX21NHSX4_S_R_Z_R 0.1
`define F_MUX21NHSX4_B_F_Z_R 0.1
`define F_MUX21NHSX4_B_R_Z_F 0.1
`define F_MUX21NHSX4_A_F_Z_R 0.1
`define F_MUX21NHSX4_A_R_Z_F 0.1

module F_MUX21NHSX4 (Z, A, B, S);

   output Z;
   input A;
   input B;
   input S;


   not  u0 (AX, A);
   not  u1 (BX, B);
   U_MUX2  u2 (Z, AX, BX, S);


   buf u3 (ST, S);
   buf u4 (BT, B);
   buf u5 (AT, A);
 
`ifdef tristatecheck
always @(ST or AT or BT)
  begin
        if (((B === 1'bz) && (S == 1)) || ((A === 1'bz) && (S == 0)) || ((S === 1'bx) && ((A === 1'bz) || (B === 1'bz))))
        $display ("WARNING: Cell F_MUX21NHSX4 used in IDDQ unsafe mode with A = %b, B = %b, S = %b at time %d", A, B, S,$time);
  end
`endif

`ifdef functional
`else
   specify

      if (!A && B) (S -=> Z) = (`F_MUX21NHSX4_S_F_Z_R,`F_MUX21NHSX4_S_R_Z_F);
      if (A && !B) (S +=> Z) = (`F_MUX21NHSX4_S_R_Z_R,`F_MUX21NHSX4_S_F_Z_F);
      (B -=> Z) = (`F_MUX21NHSX4_B_F_Z_R,`F_MUX21NHSX4_B_R_Z_F);
      (A -=> Z) = (`F_MUX21NHSX4_A_F_Z_R,`F_MUX21NHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // F_MUX21NHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:18:47 and Version :1.1 //
 
//  START 
// CELL MUX22HS 

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define MUX22HS_S_F_ZN_R 0.1
`define MUX22HS_S_R_ZN_F 0.1
`define MUX22HS_S_F_ZN_F 0.1
`define MUX22HS_S_R_ZN_R 0.1
`define MUX22HS_B_F_ZN_R 0.1
`define MUX22HS_B_R_ZN_F 0.1
`define MUX22HS_A_F_ZN_R 0.1
`define MUX22HS_A_R_ZN_F 0.1
`define MUX22HS_S_F_Z_F 0.1
`define MUX22HS_S_R_Z_R 0.1
`define MUX22HS_S_F_Z_R 0.1
`define MUX22HS_S_R_Z_F 0.1
`define MUX22HS_B_F_Z_F 0.1
`define MUX22HS_B_R_Z_R 0.1
`define MUX22HS_A_F_Z_F 0.1
`define MUX22HS_A_R_Z_R 0.1

module MUX22HS (Z, ZN, A, B, S);

   output Z;
   output ZN;
   input A;
   input B;
   input S;


   U_MUX2  u0 (Z, A, B, S);
   U_MUX2  u1 (ZN, AX, BX, S);
   not  u2 (BX, B);
   not  u3 (AX, A);

   buf u4 (ST, S);
   buf u5 (BT, B);
   buf u6 (AT, A);
 
`ifdef tristatecheck
always @(ST or AT or BT)
  begin
        if (((B === 1'bz) && (S == 1)) || ((A === 1'bz) && (S == 0)) || ((S === 1'bx) && ((A === 1'bz) || (B === 1'bz))))
        $display ("WARNING: Cell MUX22HS used in IDDQ unsafe mode with A = %b, B = %b, S = %b at time %d", A, B, S,$time);
  end
`endif

`ifdef functional
`else
   specify

      if (!A && B) (S -=> ZN) = (`MUX22HS_S_F_ZN_R,`MUX22HS_S_R_ZN_F);
      if (A && !B) (S +=> ZN) = (`MUX22HS_S_R_ZN_R,`MUX22HS_S_F_ZN_F);
      (B -=> ZN) = (`MUX22HS_B_F_ZN_R,`MUX22HS_B_R_ZN_F);
      (A -=> ZN) = (`MUX22HS_A_F_ZN_R,`MUX22HS_A_R_ZN_F);
      if (!A && B) (S +=> Z) = (`MUX22HS_S_R_Z_R,`MUX22HS_S_F_Z_F);
      if (A && !B) (S -=> Z) = (`MUX22HS_S_F_Z_R,`MUX22HS_S_R_Z_F);
      (B +=> Z) = (`MUX22HS_B_R_Z_R,`MUX22HS_B_F_Z_F);
      (A +=> Z) = (`MUX22HS_A_R_Z_R,`MUX22HS_A_F_Z_F);

   endspecify
`endif


endmodule // MUX22HS

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
//  END
// Created from CVS on Date :1998/07/07 13:19:05 and Version :1.1 //
 
//  START
// CELL MUX22HSP 

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define MUX22HSP_S_F_ZN_R 0.1
`define MUX22HSP_S_R_ZN_F 0.1
`define MUX22HSP_S_F_ZN_F 0.1
`define MUX22HSP_S_R_ZN_R 0.1
`define MUX22HSP_B_F_ZN_R 0.1
`define MUX22HSP_B_R_ZN_F 0.1
`define MUX22HSP_A_F_ZN_R 0.1
`define MUX22HSP_A_R_ZN_F 0.1
`define MUX22HSP_S_F_Z_F 0.1
`define MUX22HSP_S_R_Z_R 0.1
`define MUX22HSP_S_F_Z_R 0.1
`define MUX22HSP_S_R_Z_F 0.1
`define MUX22HSP_B_F_Z_F 0.1
`define MUX22HSP_B_R_Z_R 0.1
`define MUX22HSP_A_F_Z_F 0.1
`define MUX22HSP_A_R_Z_R 0.1

module MUX22HSP (Z, ZN, A, B, S);

   output Z;
   output ZN;
   input A;
   input B;
   input S;


   U_MUX2  u0 (Z, A, B, S);
   U_MUX2  u1 (ZN, AX, BX, S);
   not  u2 (BX, B);
   not  u3 (AX, A);

   buf u4 (ST, S);
   buf u5 (BT, B);
   buf u6 (AT, A);
 
`ifdef tristatecheck
always @(ST or AT or BT)
  begin
        if (((B === 1'bz) && (S == 1)) || ((A === 1'bz) && (S == 0)) || ((S === 1'bx) && ((A === 1'bz) || (B === 1'bz))))
        $display ("WARNING: Cell MUX22HSP used in IDDQ unsafe mode with A = %b, B = %b, S = %b at time %d", A, B, S,$time);
  end
`endif

`ifdef functional
`else
   specify

      if (!A && B) (S -=> ZN) = (`MUX22HSP_S_F_ZN_R,`MUX22HSP_S_R_ZN_F);
      if (A && !B) (S +=> ZN) = (`MUX22HSP_S_R_ZN_R,`MUX22HSP_S_F_ZN_F);
      (B -=> ZN) = (`MUX22HSP_B_F_ZN_R,`MUX22HSP_B_R_ZN_F);
      (A -=> ZN) = (`MUX22HSP_A_F_ZN_R,`MUX22HSP_A_R_ZN_F);
      if (!A && B) (S +=> Z) = (`MUX22HSP_S_R_Z_R,`MUX22HSP_S_F_Z_F);
      if (A && !B) (S -=> Z) = (`MUX22HSP_S_F_Z_R,`MUX22HSP_S_R_Z_F);
      (B +=> Z) = (`MUX22HSP_B_R_Z_R,`MUX22HSP_B_F_Z_F);
      (A +=> Z) = (`MUX22HSP_A_R_Z_R,`MUX22HSP_A_F_Z_F);

   endspecify
`endif


endmodule // MUX22HSP

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
//  END
// Created from CVS on Date :1998/07/07 13:19:05 and Version :1.1 //
 
//  START
// CELL F_MUX22HS 

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define F_MUX22HS_S_F_ZN_R 0.1
`define F_MUX22HS_S_R_ZN_F 0.1
`define F_MUX22HS_S_F_ZN_F 0.1
`define F_MUX22HS_S_R_ZN_R 0.1
`define F_MUX22HS_B_F_ZN_R 0.1
`define F_MUX22HS_B_R_ZN_F 0.1
`define F_MUX22HS_A_F_ZN_R 0.1
`define F_MUX22HS_A_R_ZN_F 0.1
`define F_MUX22HS_S_F_Z_F 0.1
`define F_MUX22HS_S_R_Z_R 0.1
`define F_MUX22HS_S_F_Z_R 0.1
`define F_MUX22HS_S_R_Z_F 0.1
`define F_MUX22HS_B_F_Z_F 0.1
`define F_MUX22HS_B_R_Z_R 0.1
`define F_MUX22HS_A_F_Z_F 0.1
`define F_MUX22HS_A_R_Z_R 0.1

module F_MUX22HS (Z, ZN, A, B, S);

   output Z;
   output ZN;
   input A;
   input B;
   input S;


   U_MUX2  u0 (Z, A, B, S);
   U_MUX2  u1 (ZN, AX, BX, S);
   not  u2 (BX, B);
   not  u3 (AX, A);

   buf u4 (ST, S);
   buf u5 (BT, B);
   buf u6 (AT, A);
 
`ifdef tristatecheck
always @(ST or AT or BT)
  begin
        if (((B === 1'bz) && (S == 1)) || ((A === 1'bz) && (S == 0)) || ((S === 1'bx) && ((A === 1'bz) || (B === 1'bz))))
        $display ("WARNING: Cell F_MUX22HS used in IDDQ unsafe mode with A = %b, B = %b, S = %b at time %d", A, B, S,$time);
  end
`endif

`ifdef functional
`else
   specify

      if (!A && B) (S -=> ZN) = (`F_MUX22HS_S_F_ZN_R,`F_MUX22HS_S_R_ZN_F);
      if (A && !B) (S +=> ZN) = (`F_MUX22HS_S_R_ZN_R,`F_MUX22HS_S_F_ZN_F);
      (B -=> ZN) = (`F_MUX22HS_B_F_ZN_R,`F_MUX22HS_B_R_ZN_F);
      (A -=> ZN) = (`F_MUX22HS_A_F_ZN_R,`F_MUX22HS_A_R_ZN_F);
      if (!A && B) (S +=> Z) = (`F_MUX22HS_S_R_Z_R,`F_MUX22HS_S_F_Z_F);
      if (A && !B) (S -=> Z) = (`F_MUX22HS_S_F_Z_R,`F_MUX22HS_S_R_Z_F);
      (B +=> Z) = (`F_MUX22HS_B_R_Z_R,`F_MUX22HS_B_F_Z_F);
      (A +=> Z) = (`F_MUX22HS_A_R_Z_R,`F_MUX22HS_A_F_Z_F);

   endspecify
`endif


endmodule // F_MUX22HS

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
//  END
// Created from CVS on Date :1998/07/07 13:19:05 and Version :1.1 //
 
//  START
// CELL F_MUX22HSP 

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define F_MUX22HSP_S_F_ZN_R 0.1
`define F_MUX22HSP_S_R_ZN_F 0.1
`define F_MUX22HSP_S_F_ZN_F 0.1
`define F_MUX22HSP_S_R_ZN_R 0.1
`define F_MUX22HSP_B_F_ZN_R 0.1
`define F_MUX22HSP_B_R_ZN_F 0.1
`define F_MUX22HSP_A_F_ZN_R 0.1
`define F_MUX22HSP_A_R_ZN_F 0.1
`define F_MUX22HSP_S_F_Z_F 0.1
`define F_MUX22HSP_S_R_Z_R 0.1
`define F_MUX22HSP_S_F_Z_R 0.1
`define F_MUX22HSP_S_R_Z_F 0.1
`define F_MUX22HSP_B_F_Z_F 0.1
`define F_MUX22HSP_B_R_Z_R 0.1
`define F_MUX22HSP_A_F_Z_F 0.1
`define F_MUX22HSP_A_R_Z_R 0.1

module F_MUX22HSP (Z, ZN, A, B, S);

   output Z;
   output ZN;
   input A;
   input B;
   input S;


   U_MUX2  u0 (Z, A, B, S);
   U_MUX2  u1 (ZN, AX, BX, S);
   not  u2 (BX, B);
   not  u3 (AX, A);

   buf u4 (ST, S);
   buf u5 (BT, B);
   buf u6 (AT, A);
 
`ifdef tristatecheck
always @(ST or AT or BT)
  begin
        if (((B === 1'bz) && (S == 1)) || ((A === 1'bz) && (S == 0)) || ((S === 1'bx) && ((A === 1'bz) || (B === 1'bz))))
        $display ("WARNING: Cell F_MUX22HSP used in IDDQ unsafe mode with A = %b, B = %b, S = %b at time %d", A, B, S,$time);
  end
`endif

`ifdef functional
`else
   specify

      if (!A && B) (S -=> ZN) = (`F_MUX22HSP_S_F_ZN_R,`F_MUX22HSP_S_R_ZN_F);
      if (A && !B) (S +=> ZN) = (`F_MUX22HSP_S_R_ZN_R,`F_MUX22HSP_S_F_ZN_F);
      (B -=> ZN) = (`F_MUX22HSP_B_F_ZN_R,`F_MUX22HSP_B_R_ZN_F);
      (A -=> ZN) = (`F_MUX22HSP_A_F_ZN_R,`F_MUX22HSP_A_R_ZN_F);
      if (!A && B) (S +=> Z) = (`F_MUX22HSP_S_R_Z_R,`F_MUX22HSP_S_F_Z_F);
      if (A && !B) (S -=> Z) = (`F_MUX22HSP_S_F_Z_R,`F_MUX22HSP_S_R_Z_F);
      (B +=> Z) = (`F_MUX22HSP_B_R_Z_R,`F_MUX22HSP_B_F_Z_F);
      (A +=> Z) = (`F_MUX22HSP_A_R_Z_R,`F_MUX22HSP_A_F_Z_F);

   endspecify
`endif


endmodule // F_MUX22HSP

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
//  END
// Created from CVS on Date :1998/07/07 13:19:05 and Version :1.1 //
 
//  START
// CELL MUX41HSX05 

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define MUX41HSX05_B_F_Z_F 0.1
`define MUX41HSX05_B_R_Z_R 0.1
`define MUX41HSX05_B_F_Z_R 0.1
`define MUX41HSX05_B_R_Z_F 0.1
`define MUX41HSX05_A_F_Z_F 0.1
`define MUX41HSX05_A_R_Z_R 0.1
`define MUX41HSX05_A_F_Z_R 0.1
`define MUX41HSX05_A_R_Z_F 0.1
`define MUX41HSX05_D3_F_Z_F 0.1
`define MUX41HSX05_D3_R_Z_R 0.1
`define MUX41HSX05_D2_F_Z_F 0.1
`define MUX41HSX05_D2_R_Z_R 0.1
`define MUX41HSX05_D1_F_Z_F 0.1
`define MUX41HSX05_D1_R_Z_R 0.1
`define MUX41HSX05_D0_F_Z_F 0.1
`define MUX41HSX05_D0_R_Z_R 0.1

module MUX41HSX05 (Z, D0, D1, D2, D3, A, B);

   output Z;
   input D0;
   input D1;
   input D2;
   input D3;
   input A;
   input B;


   // gate-level netlist replaced by UDP - 19 DEC 1995
   U_MUX4  u0 (Z, D0, D1, D2, D3, A, B);

   buf u1 (D3T, D3);
   buf u2 (D2T, D2);
   buf u3 (D1T, D1);
   buf u4 (D0T, D0);
   buf u5 (BT, B);
   buf u6 (AT, A);
 
`ifdef tristatecheck
always @(D0T or D1T or D2T or D3T or AT or BT)
begin
case ({B,A})
2'b00 : if (D0 === 1'bz)
                $display ("WARNING: Cell MUX41HSX05 used in IDDQ unsafe mode with A = %b, B = %b, D0 = %b at time %d", A, B, D0, $time);
2'b01 : if (D1 === 1'bz)
                $display ("WARNING: Cell MUX41HSX05 used in IDDQ unsafe mode with A = %b, B = %b, D1 = %b at time %d", A, B, D1, $time);
2'b10 : if (D2 === 1'bz)
                $display ("WARNING: Cell MUX41HSX05 used in IDDQ unsafe mode with A = %b, B = %b, D2 = %b at time %d", A, B, D2, $time);
2'b11 : if (D3 === 1'bz)
                $display ("WARNING: Cell MUX41HSX05 used in IDDQ unsafe mode with A = %b, B = %b, D3 = %b at time %d", A, B, D3, $time);
default:;
endcase
if (((A === 1'bx) || (B === 1'bx)) && ((D0 === 1'bz) || (D1 === 1'bz) || (D2 === 1'bz) || (D3 === 1'bz)))
begin
        $display ("WARNING: Cell MUX41HSX05 used in IDDQ unsafe mode at time %d", $time);
        $display ("         with inputs at A = %b, B = %b, D0 = %b, D1 =%b, D2 = %b, D3 = %b", A, B, D0, D1, D2, D3);
end
end
`endif
 


`ifdef functional
`else
   specify

      if (!D1 && D3 && A || !D0 && D2 && !A) (B +=> Z) = (`MUX41HSX05_B_R_Z_R,`MUX41HSX05_B_F_Z_F);
      if (D1 && !D3 && A || D0 && !D2 && !A) (B -=> Z) = (`MUX41HSX05_B_F_Z_R,`MUX41HSX05_B_R_Z_F);
      if (!D2 && D3 && B || !D0 && D1 && !B) (A +=> Z) = (`MUX41HSX05_A_R_Z_R,`MUX41HSX05_A_F_Z_F);
      if (D2 && !D3 && B || D0 && !D1 && !B) (A -=> Z) = (`MUX41HSX05_A_F_Z_R,`MUX41HSX05_A_R_Z_F);
      (D3 +=> Z) = (`MUX41HSX05_D3_R_Z_R,`MUX41HSX05_D3_F_Z_F);
      (D2 +=> Z) = (`MUX41HSX05_D2_R_Z_R,`MUX41HSX05_D2_F_Z_F);
      (D1 +=> Z) = (`MUX41HSX05_D1_R_Z_R,`MUX41HSX05_D1_F_Z_F);
      (D0 +=> Z) = (`MUX41HSX05_D0_R_Z_R,`MUX41HSX05_D0_F_Z_F);

   endspecify
`endif


endmodule // MUX41HSX05

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
//  END
// Created from CVS on Date :1998/07/07 13:19:05 and Version :1.1 //
 
//  START
// CELL MUX41HS 

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define MUX41HS_B_F_Z_F 0.1
`define MUX41HS_B_R_Z_R 0.1
`define MUX41HS_B_F_Z_R 0.1
`define MUX41HS_B_R_Z_F 0.1
`define MUX41HS_A_F_Z_F 0.1
`define MUX41HS_A_R_Z_R 0.1
`define MUX41HS_A_F_Z_R 0.1
`define MUX41HS_A_R_Z_F 0.1
`define MUX41HS_D3_F_Z_F 0.1
`define MUX41HS_D3_R_Z_R 0.1
`define MUX41HS_D2_F_Z_F 0.1
`define MUX41HS_D2_R_Z_R 0.1
`define MUX41HS_D1_F_Z_F 0.1
`define MUX41HS_D1_R_Z_R 0.1
`define MUX41HS_D0_F_Z_F 0.1
`define MUX41HS_D0_R_Z_R 0.1

module MUX41HS (Z, D0, D1, D2, D3, A, B);

   output Z;
   input D0;
   input D1;
   input D2;
   input D3;
   input A;
   input B;


   // gate-level netlist replaced by UDP - 19 DEC 1995
   U_MUX4  u0 (Z, D0, D1, D2, D3, A, B);

   buf u1 (D3T, D3);
   buf u2 (D2T, D2);
   buf u3 (D1T, D1);
   buf u4 (D0T, D0);
   buf u5 (BT, B);
   buf u6 (AT, A);
 
`ifdef tristatecheck
always @(D0T or D1T or D2T or D3T or AT or BT)
begin
case ({B,A})
2'b00 : if (D0 === 1'bz)
                $display ("WARNING: Cell MUX41HS used in IDDQ unsafe mode with A = %b, B = %b, D0 = %b at time %d", A, B, D0, $time);
2'b01 : if (D1 === 1'bz)
                $display ("WARNING: Cell MUX41HS used in IDDQ unsafe mode with A = %b, B = %b, D1 = %b at time %d", A, B, D1, $time);
2'b10 : if (D2 === 1'bz)
                $display ("WARNING: Cell MUX41HS used in IDDQ unsafe mode with A = %b, B = %b, D2 = %b at time %d", A, B, D2, $time);
2'b11 : if (D3 === 1'bz)
                $display ("WARNING: Cell MUX41HS used in IDDQ unsafe mode with A = %b, B = %b, D3 = %b at time %d", A, B, D3, $time);
default:;
endcase
if (((A === 1'bx) || (B === 1'bx)) && ((D0 === 1'bz) || (D1 === 1'bz) || (D2 === 1'bz) || (D3 === 1'bz)))
begin
        $display ("WARNING: Cell MUX41HS used in IDDQ unsafe mode at time %d", $time);
        $display ("         with inputs at A = %b, B = %b, D0 = %b, D1 =%b, D2 = %b, D3 = %b", A, B, D0, D1, D2, D3);
end
end
`endif
 


`ifdef functional
`else
   specify

      if (!D1 && D3 && A || !D0 && D2 && !A) (B +=> Z) = (`MUX41HS_B_R_Z_R,`MUX41HS_B_F_Z_F);
      if (D1 && !D3 && A || D0 && !D2 && !A) (B -=> Z) = (`MUX41HS_B_F_Z_R,`MUX41HS_B_R_Z_F);
      if (!D2 && D3 && B || !D0 && D1 && !B) (A +=> Z) = (`MUX41HS_A_R_Z_R,`MUX41HS_A_F_Z_F);
      if (D2 && !D3 && B || D0 && !D1 && !B) (A -=> Z) = (`MUX41HS_A_F_Z_R,`MUX41HS_A_R_Z_F);
      (D3 +=> Z) = (`MUX41HS_D3_R_Z_R,`MUX41HS_D3_F_Z_F);
      (D2 +=> Z) = (`MUX41HS_D2_R_Z_R,`MUX41HS_D2_F_Z_F);
      (D1 +=> Z) = (`MUX41HS_D1_R_Z_R,`MUX41HS_D1_F_Z_F);
      (D0 +=> Z) = (`MUX41HS_D0_R_Z_R,`MUX41HS_D0_F_Z_F);

   endspecify
`endif


endmodule // MUX41HS

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
//  END
// Created from CVS on Date :1998/07/07 13:19:05 and Version :1.1 //
 
//  START
// CELL MUX41HSP 

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define MUX41HSP_B_F_Z_F 0.1
`define MUX41HSP_B_R_Z_R 0.1
`define MUX41HSP_B_F_Z_R 0.1
`define MUX41HSP_B_R_Z_F 0.1
`define MUX41HSP_A_F_Z_F 0.1
`define MUX41HSP_A_R_Z_R 0.1
`define MUX41HSP_A_F_Z_R 0.1
`define MUX41HSP_A_R_Z_F 0.1
`define MUX41HSP_D3_F_Z_F 0.1
`define MUX41HSP_D3_R_Z_R 0.1
`define MUX41HSP_D2_F_Z_F 0.1
`define MUX41HSP_D2_R_Z_R 0.1
`define MUX41HSP_D1_F_Z_F 0.1
`define MUX41HSP_D1_R_Z_R 0.1
`define MUX41HSP_D0_F_Z_F 0.1
`define MUX41HSP_D0_R_Z_R 0.1

module MUX41HSP (Z, D0, D1, D2, D3, A, B);

   output Z;
   input D0;
   input D1;
   input D2;
   input D3;
   input A;
   input B;


   // gate-level netlist replaced by UDP - 19 DEC 1995
   U_MUX4  u0 (Z, D0, D1, D2, D3, A, B);

   buf u1 (D3T, D3);
   buf u2 (D2T, D2);
   buf u3 (D1T, D1);
   buf u4 (D0T, D0);
   buf u5 (BT, B);
   buf u6 (AT, A);
 
`ifdef tristatecheck
always @(D0T or D1T or D2T or D3T or AT or BT)
begin
case ({B,A})
2'b00 : if (D0 === 1'bz)
                $display ("WARNING: Cell MUX41HSP used in IDDQ unsafe mode with A = %b, B = %b, D0 = %b at time %d", A, B, D0, $time);
2'b01 : if (D1 === 1'bz)
                $display ("WARNING: Cell MUX41HSP used in IDDQ unsafe mode with A = %b, B = %b, D1 = %b at time %d", A, B, D1, $time);
2'b10 : if (D2 === 1'bz)
                $display ("WARNING: Cell MUX41HSP used in IDDQ unsafe mode with A = %b, B = %b, D2 = %b at time %d", A, B, D2, $time);
2'b11 : if (D3 === 1'bz)
                $display ("WARNING: Cell MUX41HSP used in IDDQ unsafe mode with A = %b, B = %b, D3 = %b at time %d", A, B, D3, $time);
default:;
endcase
if (((A === 1'bx) || (B === 1'bx)) && ((D0 === 1'bz) || (D1 === 1'bz) || (D2 === 1'bz) || (D3 === 1'bz)))
begin
        $display ("WARNING: Cell MUX41HSP used in IDDQ unsafe mode at time %d", $time);
        $display ("         with inputs at A = %b, B = %b, D0 = %b, D1 =%b, D2 = %b, D3 = %b", A, B, D0, D1, D2, D3);
end
end
`endif
 


`ifdef functional
`else
   specify

      if (!D1 && D3 && A || !D0 && D2 && !A) (B +=> Z) = (`MUX41HSP_B_R_Z_R,`MUX41HSP_B_F_Z_F);
      if (D1 && !D3 && A || D0 && !D2 && !A) (B -=> Z) = (`MUX41HSP_B_F_Z_R,`MUX41HSP_B_R_Z_F);
      if (!D2 && D3 && B || !D0 && D1 && !B) (A +=> Z) = (`MUX41HSP_A_R_Z_R,`MUX41HSP_A_F_Z_F);
      if (D2 && !D3 && B || D0 && !D1 && !B) (A -=> Z) = (`MUX41HSP_A_F_Z_R,`MUX41HSP_A_R_Z_F);
      (D3 +=> Z) = (`MUX41HSP_D3_R_Z_R,`MUX41HSP_D3_F_Z_F);
      (D2 +=> Z) = (`MUX41HSP_D2_R_Z_R,`MUX41HSP_D2_F_Z_F);
      (D1 +=> Z) = (`MUX41HSP_D1_R_Z_R,`MUX41HSP_D1_F_Z_F);
      (D0 +=> Z) = (`MUX41HSP_D0_R_Z_R,`MUX41HSP_D0_F_Z_F);

   endspecify
`endif


endmodule // MUX41HSP

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
//  END
// Created from CVS on Date :1998/07/07 13:19:05 and Version :1.1 //
 
//  START
// CELL MUX41HSX4 

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define MUX41HSX4_B_F_Z_F 0.1
`define MUX41HSX4_B_R_Z_R 0.1
`define MUX41HSX4_B_F_Z_R 0.1
`define MUX41HSX4_B_R_Z_F 0.1
`define MUX41HSX4_A_F_Z_F 0.1
`define MUX41HSX4_A_R_Z_R 0.1
`define MUX41HSX4_A_F_Z_R 0.1
`define MUX41HSX4_A_R_Z_F 0.1
`define MUX41HSX4_D3_F_Z_F 0.1
`define MUX41HSX4_D3_R_Z_R 0.1
`define MUX41HSX4_D2_F_Z_F 0.1
`define MUX41HSX4_D2_R_Z_R 0.1
`define MUX41HSX4_D1_F_Z_F 0.1
`define MUX41HSX4_D1_R_Z_R 0.1
`define MUX41HSX4_D0_F_Z_F 0.1
`define MUX41HSX4_D0_R_Z_R 0.1

module MUX41HSX4 (Z, D0, D1, D2, D3, A, B);

   output Z;
   input D0;
   input D1;
   input D2;
   input D3;
   input A;
   input B;


   // gate-level netlist replaced by UDP - 19 DEC 1995
   U_MUX4  u0 (Z, D0, D1, D2, D3, A, B);

   buf u1 (D3T, D3);
   buf u2 (D2T, D2);
   buf u3 (D1T, D1);
   buf u4 (D0T, D0);
   buf u5 (BT, B);
   buf u6 (AT, A);
 
`ifdef tristatecheck
always @(D0T or D1T or D2T or D3T or AT or BT)
begin
case ({B,A})
2'b00 : if (D0 === 1'bz)
                $display ("WARNING: Cell MUX41HSX4 used in IDDQ unsafe mode with A = %b, B = %b, D0 = %b at time %d", A, B, D0, $time);
2'b01 : if (D1 === 1'bz)
                $display ("WARNING: Cell MUX41HSX4 used in IDDQ unsafe mode with A = %b, B = %b, D1 = %b at time %d", A, B, D1, $time);
2'b10 : if (D2 === 1'bz)
                $display ("WARNING: Cell MUX41HSX4 used in IDDQ unsafe mode with A = %b, B = %b, D2 = %b at time %d", A, B, D2, $time);
2'b11 : if (D3 === 1'bz)
                $display ("WARNING: Cell MUX41HSX4 used in IDDQ unsafe mode with A = %b, B = %b, D3 = %b at time %d", A, B, D3, $time);
default:;
endcase
if (((A === 1'bx) || (B === 1'bx)) && ((D0 === 1'bz) || (D1 === 1'bz) || (D2 === 1'bz) || (D3 === 1'bz)))
begin
        $display ("WARNING: Cell MUX41HSX4 used in IDDQ unsafe mode at time %d", $time);
        $display ("         with inputs at A = %b, B = %b, D0 = %b, D1 =%b, D2 = %b, D3 = %b", A, B, D0, D1, D2, D3);
end
end
`endif
 


`ifdef functional
`else
   specify

      if (!D1 && D3 && A || !D0 && D2 && !A) (B +=> Z) = (`MUX41HSX4_B_R_Z_R,`MUX41HSX4_B_F_Z_F);
      if (D1 && !D3 && A || D0 && !D2 && !A) (B -=> Z) = (`MUX41HSX4_B_F_Z_R,`MUX41HSX4_B_R_Z_F);
      if (!D2 && D3 && B || !D0 && D1 && !B) (A +=> Z) = (`MUX41HSX4_A_R_Z_R,`MUX41HSX4_A_F_Z_F);
      if (D2 && !D3 && B || D0 && !D1 && !B) (A -=> Z) = (`MUX41HSX4_A_F_Z_R,`MUX41HSX4_A_R_Z_F);
      (D3 +=> Z) = (`MUX41HSX4_D3_R_Z_R,`MUX41HSX4_D3_F_Z_F);
      (D2 +=> Z) = (`MUX41HSX4_D2_R_Z_R,`MUX41HSX4_D2_F_Z_F);
      (D1 +=> Z) = (`MUX41HSX4_D1_R_Z_R,`MUX41HSX4_D1_F_Z_F);
      (D0 +=> Z) = (`MUX41HSX4_D0_R_Z_R,`MUX41HSX4_D0_F_Z_F);

   endspecify
`endif


endmodule // MUX41HSX4

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
//  END
// Created from CVS on Date :1998/07/07 13:19:05 and Version :1.1 //
 
//  START
// CELL MUX41NHS 

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define MUX41NHS_B_F_Z_R 0.1
`define MUX41NHS_B_R_Z_F 0.1
`define MUX41NHS_B_F_Z_F 0.1
`define MUX41NHS_B_R_Z_R 0.1
`define MUX41NHS_A_F_Z_R 0.1
`define MUX41NHS_A_R_Z_F 0.1
`define MUX41NHS_A_F_Z_F 0.1
`define MUX41NHS_A_R_Z_R 0.1
`define MUX41NHS_D3_F_Z_R 0.1
`define MUX41NHS_D3_R_Z_F 0.1
`define MUX41NHS_D2_F_Z_R 0.1
`define MUX41NHS_D2_R_Z_F 0.1
`define MUX41NHS_D1_F_Z_R 0.1
`define MUX41NHS_D1_R_Z_F 0.1
`define MUX41NHS_D0_F_Z_R 0.1
`define MUX41NHS_D0_R_Z_F 0.1

module MUX41NHS (Z, D0, D1, D2, D3, A, B);

   output Z;
   input D0;
   input D1;
   input D2;
   input D3;
   input A;
   input B;


   // gate-level netlist replaced by UDP - 19 DEC 1995
   U_MUX4  u0 (ZX, D0, D1, D2, D3, A, B);
   not  u7 (Z, ZX);

   buf u1 (D3T, D3);
   buf u2 (D2T, D2);
   buf u3 (D1T, D1);
   buf u4 (D0T, D0);
   buf u5 (BT, B);
   buf u6 (AT, A);
 
`ifdef tristatecheck
always @(D0T or D1T or D2T or D3T or AT or BT)
begin
case ({B,A})
2'b00 : if (D0 === 1'bz)
                $display ("WARNING: Cell MUX41NHS used in IDDQ unsafe mode with A = %b, B = %b, D0 = %b at time %d", A, B, D0, $time);
2'b01 : if (D1 === 1'bz)
                $display ("WARNING: Cell MUX41NHS used in IDDQ unsafe mode with A = %b, B = %b, D1 = %b at time %d", A, B, D1, $time);
2'b10 : if (D2 === 1'bz)
                $display ("WARNING: Cell MUX41NHS used in IDDQ unsafe mode with A = %b, B = %b, D2 = %b at time %d", A, B, D2, $time);
2'b11 : if (D3 === 1'bz)
                $display ("WARNING: Cell MUX41NHS used in IDDQ unsafe mode with A = %b, B = %b, D3 = %b at time %d", A, B, D3, $time);
default:;
endcase
if (((A === 1'bx) || (B === 1'bx)) && ((D0 === 1'bz) || (D1 === 1'bz) || (D2 === 1'bz) || (D3 === 1'bz)))
begin
        $display ("WARNING: Cell MUX41NHS used in IDDQ unsafe mode at time %d", $time);
        $display ("         with inputs at A = %b, B = %b, D0 = %b, D1 =%b, D2 = %b, D3 = %b", A, B, D0, D1, D2, D3);
end
end
`endif
 


`ifdef functional
`else
   specify

      if (!D1 && D3 && A || !D0 && D2 && !A) (B -=> Z) = (`MUX41NHS_B_F_Z_R,`MUX41NHS_B_R_Z_F);
      if (D1 && !D3 && A || D0 && !D2 && !A) (B +=> Z) = (`MUX41NHS_B_R_Z_R,`MUX41NHS_B_F_Z_F);
      if (!D2 && D3 && B || !D0 && D1 && !B) (A -=> Z) = (`MUX41NHS_A_F_Z_R,`MUX41NHS_A_R_Z_F);
      if (D2 && !D3 && B || D0 && !D1 && !B) (A +=> Z) = (`MUX41NHS_A_R_Z_R,`MUX41NHS_A_F_Z_F);
      (D3 -=> Z) = (`MUX41NHS_D3_F_Z_R,`MUX41NHS_D3_R_Z_F);
      (D2 -=> Z) = (`MUX41NHS_D2_F_Z_R,`MUX41NHS_D2_R_Z_F);
      (D1 -=> Z) = (`MUX41NHS_D1_F_Z_R,`MUX41NHS_D1_R_Z_F);
      (D0 -=> Z) = (`MUX41NHS_D0_F_Z_R,`MUX41NHS_D0_R_Z_F);

   endspecify
`endif


endmodule // MUX41NHS

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
//  END
// Created from CVS on Date :1998/07/07 13:19:05 and Version :1.1 //
 
//  START
// CELL MUX41NHSP 

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define MUX41NHSP_B_F_Z_R 0.1
`define MUX41NHSP_B_R_Z_F 0.1
`define MUX41NHSP_B_F_Z_F 0.1
`define MUX41NHSP_B_R_Z_R 0.1
`define MUX41NHSP_A_F_Z_R 0.1
`define MUX41NHSP_A_R_Z_F 0.1
`define MUX41NHSP_A_F_Z_F 0.1
`define MUX41NHSP_A_R_Z_R 0.1
`define MUX41NHSP_D3_F_Z_R 0.1
`define MUX41NHSP_D3_R_Z_F 0.1
`define MUX41NHSP_D2_F_Z_R 0.1
`define MUX41NHSP_D2_R_Z_F 0.1
`define MUX41NHSP_D1_F_Z_R 0.1
`define MUX41NHSP_D1_R_Z_F 0.1
`define MUX41NHSP_D0_F_Z_R 0.1
`define MUX41NHSP_D0_R_Z_F 0.1

module MUX41NHSP (Z, D0, D1, D2, D3, A, B);

   output Z;
   input D0;
   input D1;
   input D2;
   input D3;
   input A;
   input B;


   // gate-level netlist replaced by UDP - 19 DEC 1995
   U_MUX4  u0 (ZX, D0, D1, D2, D3, A, B);
   not  u7 (Z, ZX);

   buf u1 (D3T, D3);
   buf u2 (D2T, D2);
   buf u3 (D1T, D1);
   buf u4 (D0T, D0);
   buf u5 (BT, B);
   buf u6 (AT, A);
 
`ifdef tristatecheck
always @(D0T or D1T or D2T or D3T or AT or BT)
begin
case ({B,A})
2'b00 : if (D0 === 1'bz)
                $display ("WARNING: Cell MUX41NHSP used in IDDQ unsafe mode with A = %b, B = %b, D0 = %b at time %d", A, B, D0, $time);
2'b01 : if (D1 === 1'bz)
                $display ("WARNING: Cell MUX41NHSP used in IDDQ unsafe mode with A = %b, B = %b, D1 = %b at time %d", A, B, D1, $time);
2'b10 : if (D2 === 1'bz)
                $display ("WARNING: Cell MUX41NHSP used in IDDQ unsafe mode with A = %b, B = %b, D2 = %b at time %d", A, B, D2, $time);
2'b11 : if (D3 === 1'bz)
                $display ("WARNING: Cell MUX41NHSP used in IDDQ unsafe mode with A = %b, B = %b, D3 = %b at time %d", A, B, D3, $time);
default:;
endcase
if (((A === 1'bx) || (B === 1'bx)) && ((D0 === 1'bz) || (D1 === 1'bz) || (D2 === 1'bz) || (D3 === 1'bz)))
begin
        $display ("WARNING: Cell MUX41NHSP used in IDDQ unsafe mode at time %d", $time);
        $display ("         with inputs at A = %b, B = %b, D0 = %b, D1 =%b, D2 = %b, D3 = %b", A, B, D0, D1, D2, D3);
end
end
`endif
 


`ifdef functional
`else
   specify

      if (!D1 && D3 && A || !D0 && D2 && !A) (B -=> Z) = (`MUX41NHSP_B_F_Z_R,`MUX41NHSP_B_R_Z_F);
      if (D1 && !D3 && A || D0 && !D2 && !A) (B +=> Z) = (`MUX41NHSP_B_R_Z_R,`MUX41NHSP_B_F_Z_F);
      if (!D2 && D3 && B || !D0 && D1 && !B) (A -=> Z) = (`MUX41NHSP_A_F_Z_R,`MUX41NHSP_A_R_Z_F);
      if (D2 && !D3 && B || D0 && !D1 && !B) (A +=> Z) = (`MUX41NHSP_A_R_Z_R,`MUX41NHSP_A_F_Z_F);
      (D3 -=> Z) = (`MUX41NHSP_D3_F_Z_R,`MUX41NHSP_D3_R_Z_F);
      (D2 -=> Z) = (`MUX41NHSP_D2_F_Z_R,`MUX41NHSP_D2_R_Z_F);
      (D1 -=> Z) = (`MUX41NHSP_D1_F_Z_R,`MUX41NHSP_D1_R_Z_F);
      (D0 -=> Z) = (`MUX41NHSP_D0_F_Z_R,`MUX41NHSP_D0_R_Z_F);

   endspecify
`endif


endmodule // MUX41NHSP

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
//  END
// Created from CVS on Date :1998/07/07 13:19:05 and Version :1.1 //
 
//  START
// CELL MUX41NHSX4 

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define MUX41NHSX4_B_F_Z_R 0.1
`define MUX41NHSX4_B_R_Z_F 0.1
`define MUX41NHSX4_B_F_Z_F 0.1
`define MUX41NHSX4_B_R_Z_R 0.1
`define MUX41NHSX4_A_F_Z_R 0.1
`define MUX41NHSX4_A_R_Z_F 0.1
`define MUX41NHSX4_A_F_Z_F 0.1
`define MUX41NHSX4_A_R_Z_R 0.1
`define MUX41NHSX4_D3_F_Z_R 0.1
`define MUX41NHSX4_D3_R_Z_F 0.1
`define MUX41NHSX4_D2_F_Z_R 0.1
`define MUX41NHSX4_D2_R_Z_F 0.1
`define MUX41NHSX4_D1_F_Z_R 0.1
`define MUX41NHSX4_D1_R_Z_F 0.1
`define MUX41NHSX4_D0_F_Z_R 0.1
`define MUX41NHSX4_D0_R_Z_F 0.1

module MUX41NHSX4 (Z, D0, D1, D2, D3, A, B);

   output Z;
   input D0;
   input D1;
   input D2;
   input D3;
   input A;
   input B;


   // gate-level netlist replaced by UDP - 19 DEC 1995
   U_MUX4  u0 (ZX, D0, D1, D2, D3, A, B);
   not  u7 (Z, ZX);

   buf u1 (D3T, D3);
   buf u2 (D2T, D2);
   buf u3 (D1T, D1);
   buf u4 (D0T, D0);
   buf u5 (BT, B);
   buf u6 (AT, A);
 
`ifdef tristatecheck
always @(D0T or D1T or D2T or D3T or AT or BT)
begin
case ({B,A})
2'b00 : if (D0 === 1'bz)
                $display ("WARNING: Cell MUX41NHSX4 used in IDDQ unsafe mode with A = %b, B = %b, D0 = %b at time %d", A, B, D0, $time);
2'b01 : if (D1 === 1'bz)
                $display ("WARNING: Cell MUX41NHSX4 used in IDDQ unsafe mode with A = %b, B = %b, D1 = %b at time %d", A, B, D1, $time);
2'b10 : if (D2 === 1'bz)
                $display ("WARNING: Cell MUX41NHSX4 used in IDDQ unsafe mode with A = %b, B = %b, D2 = %b at time %d", A, B, D2, $time);
2'b11 : if (D3 === 1'bz)
                $display ("WARNING: Cell MUX41NHSX4 used in IDDQ unsafe mode with A = %b, B = %b, D3 = %b at time %d", A, B, D3, $time);
default:;
endcase
if (((A === 1'bx) || (B === 1'bx)) && ((D0 === 1'bz) || (D1 === 1'bz) || (D2 === 1'bz) || (D3 === 1'bz)))
begin
        $display ("WARNING: Cell MUX41NHSX4 used in IDDQ unsafe mode at time %d", $time);
        $display ("         with inputs at A = %b, B = %b, D0 = %b, D1 =%b, D2 = %b, D3 = %b", A, B, D0, D1, D2, D3);
end
end
`endif
 


`ifdef functional
`else
   specify

      if (!D1 && D3 && A || !D0 && D2 && !A) (B -=> Z) = (`MUX41NHSX4_B_F_Z_R,`MUX41NHSX4_B_R_Z_F);
      if (D1 && !D3 && A || D0 && !D2 && !A) (B +=> Z) = (`MUX41NHSX4_B_R_Z_R,`MUX41NHSX4_B_F_Z_F);
      if (!D2 && D3 && B || !D0 && D1 && !B) (A -=> Z) = (`MUX41NHSX4_A_F_Z_R,`MUX41NHSX4_A_R_Z_F);
      if (D2 && !D3 && B || D0 && !D1 && !B) (A +=> Z) = (`MUX41NHSX4_A_R_Z_R,`MUX41NHSX4_A_F_Z_F);
      (D3 -=> Z) = (`MUX41NHSX4_D3_F_Z_R,`MUX41NHSX4_D3_R_Z_F);
      (D2 -=> Z) = (`MUX41NHSX4_D2_F_Z_R,`MUX41NHSX4_D2_R_Z_F);
      (D1 -=> Z) = (`MUX41NHSX4_D1_F_Z_R,`MUX41NHSX4_D1_R_Z_F);
      (D0 -=> Z) = (`MUX41NHSX4_D0_F_Z_R,`MUX41NHSX4_D0_R_Z_F);

   endspecify
`endif


endmodule // MUX41NHSX4

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
//  END
// Created from CVS on Date :1998/07/07 13:19:05 and Version :1.1 //
 
//  START
// CELL MUX81HSX05 

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define MUX81HSX05_C_F_Z_F 0.1
`define MUX81HSX05_C_R_Z_R 0.1
`define MUX81HSX05_C_F_Z_R 0.1
`define MUX81HSX05_C_R_Z_F 0.1
`define MUX81HSX05_B_F_Z_F 0.1
`define MUX81HSX05_B_R_Z_R 0.1
`define MUX81HSX05_B_F_Z_R 0.1
`define MUX81HSX05_B_R_Z_F 0.1
`define MUX81HSX05_A_F_Z_F 0.1
`define MUX81HSX05_A_R_Z_R 0.1
`define MUX81HSX05_A_F_Z_R 0.1
`define MUX81HSX05_A_R_Z_F 0.1
`define MUX81HSX05_D7_F_Z_F 0.1
`define MUX81HSX05_D7_R_Z_R 0.1
`define MUX81HSX05_D6_F_Z_F 0.1
`define MUX81HSX05_D6_R_Z_R 0.1
`define MUX81HSX05_D5_F_Z_F 0.1
`define MUX81HSX05_D5_R_Z_R 0.1
`define MUX81HSX05_D4_F_Z_F 0.1
`define MUX81HSX05_D4_R_Z_R 0.1
`define MUX81HSX05_D3_F_Z_F 0.1
`define MUX81HSX05_D3_R_Z_R 0.1
`define MUX81HSX05_D2_F_Z_F 0.1
`define MUX81HSX05_D2_R_Z_R 0.1
`define MUX81HSX05_D1_F_Z_F 0.1
`define MUX81HSX05_D1_R_Z_R 0.1
`define MUX81HSX05_D0_F_Z_F 0.1
`define MUX81HSX05_D0_R_Z_R 0.1

module MUX81HSX05 (Z, D0, D1, D2, D3, D4, D5, D6, D7, A, B, C);

   output Z;
   input D0;
   input D1;
   input D2;
   input D3;
   input D4;
   input D5;
   input D6;
   input D7;
   input A;
   input B;
   input C;


   // gate-level netlist replaced by UDPs - 19 DEC 1995
   U_MUX4    u0 (OUT_UDP_D0_TO_3_IN, D0, D1, D2, D3, A, B);
   U_MUX4    u1 (OUT_UDP_D4_TO_7_IN, D4, D5, D6, D7, A, B);
   U_MUX2  u2 (Z, OUT_UDP_D0_TO_3_IN, OUT_UDP_D4_TO_7_IN, C);

   buf u3 (D7T, D7);
   buf u4 (D6T, D6);
   buf u5 (D5T, D5);
   buf u6 (D4T, D4);
   buf u7 (D3T, D3);
   buf u8 (D2T, D2);
   buf u9 (D1T, D1);
   buf u10 (D0T, D0);
   buf u11 (CT, C);
   buf u12 (BT, B);
   buf u13 (AT, A);
 
`ifdef tristatecheck
always @(D0T or D1T or D2T or D3T or D4T or D5T or D6T or D7T or AT or BT or CT)
begin
case ({C,B,A})
3'b000 : if (D0 === 1'bz)
                $display ("WARNING: Cell MUX81HSX05 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D0 = %b at time %d", A, B, C, D0, $time);
3'b001 : if (D1 === 1'bz)
                $display ("WARNING: Cell MUX81HSX05 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D1 = %b at time %d", A, B, C, D1, $time);
3'b010 : if (D2 === 1'bz)
                $display ("WARNING: Cell MUX81HSX05 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D2 = %b at time %d", A, B, C, D2, $time);
3'b011 : if (D3 === 1'bz)
                $display ("WARNING: Cell MUX81HSX05 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D3 = %b at time %d", A, B, C, D3, $time);
3'b100 : if (D4 === 1'bz)
                $display ("WARNING: Cell MUX81HSX05 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D4 = %b at time %d", A, B, C, D4, $time);
3'b101 : if (D5 === 1'bz)
                $display ("WARNING: Cell MUX81HSX05 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D5 = %b at time %d", A, B, C, D5, $time);
3'b110 : if (D6 === 1'bz)
                $display ("WARNING: Cell MUX81HSX05 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D6 = %b at time %d", A, B, C, D6, $time);
3'b111 : if (D7 === 1'bz)
                $display ("WARNING: Cell MUX81HSX05 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D7 = %b at time %d", A, B, C, D7, $time);
default:;
endcase
if (((A === 1'bx) || (B === 1'bx) || (C === 1'bx)) && 
    ((D0 === 1'bz) || (D1 === 1'bz) || (D2 === 1'bz) || (D3 === 1'bz) || (D4 === 1'bz) || (D5 === 1'bz) || (D6 === 1'bz) || (D7 === 1'bz)))
begin
        $display ("WARNING: Cell MUX81HSX05 used in IDDQ unsafe mode at time %d", $time);
        $display ("         with inputs at A = %b, B = %b, C = %b, D0 = %b, D1 = %b, D2 = %b, D3 = %b, D4 = %b, D5 = %b, D6 = %b, D7 = %b", 
           A, B, C, D0, D1, D2, D3, D4, D5, D6, D7);
end
end
`endif


`ifdef functional
`else
   specify

      if (!D3 && D7 && A && B || !D2 && D6 && !A && B || !D1 && D5 && A && !B || !D0 && D4 && !A && !B) (C +=> Z) = (`MUX81HSX05_C_R_Z_R,`MUX81HSX05_C_F_Z_F);
      if (D3 && !D7 && A && B || D2 && !D6 && !A && B || D1 && !D5 && A && !B || D0 && !D4 && !A && !B) (C -=> Z) = (`MUX81HSX05_C_F_Z_R,`MUX81HSX05_C_R_Z_F);
      if (!D5 && D7 && A && C || !D4 && D6 && !A && C || !D1 && D3 && A && !C || !D0 && D2 && !A && !C) (B +=> Z) = (`MUX81HSX05_B_R_Z_R,`MUX81HSX05_B_F_Z_F);
      if (D5 && !D7 && A && C || D4 && !D6 && !A && C || D1 && !D3 && A && !C || D0 && !D2 && !A && !C) (B -=> Z) = (`MUX81HSX05_B_F_Z_R,`MUX81HSX05_B_R_Z_F);
      if (!D6 && D7 && B && C || !D4 && D5 && !B && C || !D2 && D3 && B && !C || !D0 && D1 && !B && !C) (A +=> Z) = (`MUX81HSX05_A_R_Z_R,`MUX81HSX05_A_F_Z_F);
      if (D6 && !D7 && B && C || D4 && !D5 && !B && C || D2 && !D3 && B && !C || D0 && !D1 && !B && !C) (A -=> Z) = (`MUX81HSX05_A_F_Z_R,`MUX81HSX05_A_R_Z_F);
      (D7 +=> Z) = (`MUX81HSX05_D7_R_Z_R,`MUX81HSX05_D7_F_Z_F);
      (D6 +=> Z) = (`MUX81HSX05_D6_R_Z_R,`MUX81HSX05_D6_F_Z_F);
      (D5 +=> Z) = (`MUX81HSX05_D5_R_Z_R,`MUX81HSX05_D5_F_Z_F);
      (D4 +=> Z) = (`MUX81HSX05_D4_R_Z_R,`MUX81HSX05_D4_F_Z_F);
      (D3 +=> Z) = (`MUX81HSX05_D3_R_Z_R,`MUX81HSX05_D3_F_Z_F);
      (D2 +=> Z) = (`MUX81HSX05_D2_R_Z_R,`MUX81HSX05_D2_F_Z_F);
      (D1 +=> Z) = (`MUX81HSX05_D1_R_Z_R,`MUX81HSX05_D1_F_Z_F);
      (D0 +=> Z) = (`MUX81HSX05_D0_R_Z_R,`MUX81HSX05_D0_F_Z_F);

   endspecify
`endif


endmodule // MUX81HSX05

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
  
//  END
// Created from CVS on Date :1998/07/07 13:19:11 and Version :1.1 //
 
//  START
// CELL MUX81HS 

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define MUX81HS_C_F_Z_F 0.1
`define MUX81HS_C_R_Z_R 0.1
`define MUX81HS_C_F_Z_R 0.1
`define MUX81HS_C_R_Z_F 0.1
`define MUX81HS_B_F_Z_F 0.1
`define MUX81HS_B_R_Z_R 0.1
`define MUX81HS_B_F_Z_R 0.1
`define MUX81HS_B_R_Z_F 0.1
`define MUX81HS_A_F_Z_F 0.1
`define MUX81HS_A_R_Z_R 0.1
`define MUX81HS_A_F_Z_R 0.1
`define MUX81HS_A_R_Z_F 0.1
`define MUX81HS_D7_F_Z_F 0.1
`define MUX81HS_D7_R_Z_R 0.1
`define MUX81HS_D6_F_Z_F 0.1
`define MUX81HS_D6_R_Z_R 0.1
`define MUX81HS_D5_F_Z_F 0.1
`define MUX81HS_D5_R_Z_R 0.1
`define MUX81HS_D4_F_Z_F 0.1
`define MUX81HS_D4_R_Z_R 0.1
`define MUX81HS_D3_F_Z_F 0.1
`define MUX81HS_D3_R_Z_R 0.1
`define MUX81HS_D2_F_Z_F 0.1
`define MUX81HS_D2_R_Z_R 0.1
`define MUX81HS_D1_F_Z_F 0.1
`define MUX81HS_D1_R_Z_R 0.1
`define MUX81HS_D0_F_Z_F 0.1
`define MUX81HS_D0_R_Z_R 0.1

module MUX81HS (Z, D0, D1, D2, D3, D4, D5, D6, D7, A, B, C);

   output Z;
   input D0;
   input D1;
   input D2;
   input D3;
   input D4;
   input D5;
   input D6;
   input D7;
   input A;
   input B;
   input C;


   // gate-level netlist replaced by UDPs - 19 DEC 1995
   U_MUX4    u0 (OUT_UDP_D0_TO_3_IN, D0, D1, D2, D3, A, B);
   U_MUX4    u1 (OUT_UDP_D4_TO_7_IN, D4, D5, D6, D7, A, B);
   U_MUX2  u2 (Z, OUT_UDP_D0_TO_3_IN, OUT_UDP_D4_TO_7_IN, C);

   buf u3 (D7T, D7);
   buf u4 (D6T, D6);
   buf u5 (D5T, D5);
   buf u6 (D4T, D4);
   buf u7 (D3T, D3);
   buf u8 (D2T, D2);
   buf u9 (D1T, D1);
   buf u10 (D0T, D0);
   buf u11 (CT, C);
   buf u12 (BT, B);
   buf u13 (AT, A);
 
`ifdef tristatecheck
always @(D0T or D1T or D2T or D3T or D4T or D5T or D6T or D7T or AT or BT or CT)
begin
case ({C,B,A})
3'b000 : if (D0 === 1'bz)
                $display ("WARNING: Cell MUX81HS used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D0 = %b at time %d", A, B, C, D0, $time);
3'b001 : if (D1 === 1'bz)
                $display ("WARNING: Cell MUX81HS used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D1 = %b at time %d", A, B, C, D1, $time);
3'b010 : if (D2 === 1'bz)
                $display ("WARNING: Cell MUX81HS used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D2 = %b at time %d", A, B, C, D2, $time);
3'b011 : if (D3 === 1'bz)
                $display ("WARNING: Cell MUX81HS used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D3 = %b at time %d", A, B, C, D3, $time);
3'b100 : if (D4 === 1'bz)
                $display ("WARNING: Cell MUX81HS used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D4 = %b at time %d", A, B, C, D4, $time);
3'b101 : if (D5 === 1'bz)
                $display ("WARNING: Cell MUX81HS used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D5 = %b at time %d", A, B, C, D5, $time);
3'b110 : if (D6 === 1'bz)
                $display ("WARNING: Cell MUX81HS used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D6 = %b at time %d", A, B, C, D6, $time);
3'b111 : if (D7 === 1'bz)
                $display ("WARNING: Cell MUX81HS used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D7 = %b at time %d", A, B, C, D7, $time);
default:;
endcase
if (((A === 1'bx) || (B === 1'bx) || (C === 1'bx)) && 
    ((D0 === 1'bz) || (D1 === 1'bz) || (D2 === 1'bz) || (D3 === 1'bz) || (D4 === 1'bz) || (D5 === 1'bz) || (D6 === 1'bz) || (D7 === 1'bz)))
begin
        $display ("WARNING: Cell MUX81HS used in IDDQ unsafe mode at time %d", $time);
        $display ("         with inputs at A = %b, B = %b, C = %b, D0 = %b, D1 = %b, D2 = %b, D3 = %b, D4 = %b, D5 = %b, D6 = %b, D7 = %b", 
           A, B, C, D0, D1, D2, D3, D4, D5, D6, D7);
end
end
`endif


`ifdef functional
`else
   specify

      if (!D3 && D7 && A && B || !D2 && D6 && !A && B || !D1 && D5 && A && !B || !D0 && D4 && !A && !B) (C +=> Z) = (`MUX81HS_C_R_Z_R,`MUX81HS_C_F_Z_F);
      if (D3 && !D7 && A && B || D2 && !D6 && !A && B || D1 && !D5 && A && !B || D0 && !D4 && !A && !B) (C -=> Z) = (`MUX81HS_C_F_Z_R,`MUX81HS_C_R_Z_F);
      if (!D5 && D7 && A && C || !D4 && D6 && !A && C || !D1 && D3 && A && !C || !D0 && D2 && !A && !C) (B +=> Z) = (`MUX81HS_B_R_Z_R,`MUX81HS_B_F_Z_F);
      if (D5 && !D7 && A && C || D4 && !D6 && !A && C || D1 && !D3 && A && !C || D0 && !D2 && !A && !C) (B -=> Z) = (`MUX81HS_B_F_Z_R,`MUX81HS_B_R_Z_F);
      if (!D6 && D7 && B && C || !D4 && D5 && !B && C || !D2 && D3 && B && !C || !D0 && D1 && !B && !C) (A +=> Z) = (`MUX81HS_A_R_Z_R,`MUX81HS_A_F_Z_F);
      if (D6 && !D7 && B && C || D4 && !D5 && !B && C || D2 && !D3 && B && !C || D0 && !D1 && !B && !C) (A -=> Z) = (`MUX81HS_A_F_Z_R,`MUX81HS_A_R_Z_F);
      (D7 +=> Z) = (`MUX81HS_D7_R_Z_R,`MUX81HS_D7_F_Z_F);
      (D6 +=> Z) = (`MUX81HS_D6_R_Z_R,`MUX81HS_D6_F_Z_F);
      (D5 +=> Z) = (`MUX81HS_D5_R_Z_R,`MUX81HS_D5_F_Z_F);
      (D4 +=> Z) = (`MUX81HS_D4_R_Z_R,`MUX81HS_D4_F_Z_F);
      (D3 +=> Z) = (`MUX81HS_D3_R_Z_R,`MUX81HS_D3_F_Z_F);
      (D2 +=> Z) = (`MUX81HS_D2_R_Z_R,`MUX81HS_D2_F_Z_F);
      (D1 +=> Z) = (`MUX81HS_D1_R_Z_R,`MUX81HS_D1_F_Z_F);
      (D0 +=> Z) = (`MUX81HS_D0_R_Z_R,`MUX81HS_D0_F_Z_F);

   endspecify
`endif


endmodule // MUX81HS

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
  
//  END
// Created from CVS on Date :1998/07/07 13:19:11 and Version :1.1 //
 
//  START
// CELL MUX81HSP 

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define MUX81HSP_C_F_Z_F 0.1
`define MUX81HSP_C_R_Z_R 0.1
`define MUX81HSP_C_F_Z_R 0.1
`define MUX81HSP_C_R_Z_F 0.1
`define MUX81HSP_B_F_Z_F 0.1
`define MUX81HSP_B_R_Z_R 0.1
`define MUX81HSP_B_F_Z_R 0.1
`define MUX81HSP_B_R_Z_F 0.1
`define MUX81HSP_A_F_Z_F 0.1
`define MUX81HSP_A_R_Z_R 0.1
`define MUX81HSP_A_F_Z_R 0.1
`define MUX81HSP_A_R_Z_F 0.1
`define MUX81HSP_D7_F_Z_F 0.1
`define MUX81HSP_D7_R_Z_R 0.1
`define MUX81HSP_D6_F_Z_F 0.1
`define MUX81HSP_D6_R_Z_R 0.1
`define MUX81HSP_D5_F_Z_F 0.1
`define MUX81HSP_D5_R_Z_R 0.1
`define MUX81HSP_D4_F_Z_F 0.1
`define MUX81HSP_D4_R_Z_R 0.1
`define MUX81HSP_D3_F_Z_F 0.1
`define MUX81HSP_D3_R_Z_R 0.1
`define MUX81HSP_D2_F_Z_F 0.1
`define MUX81HSP_D2_R_Z_R 0.1
`define MUX81HSP_D1_F_Z_F 0.1
`define MUX81HSP_D1_R_Z_R 0.1
`define MUX81HSP_D0_F_Z_F 0.1
`define MUX81HSP_D0_R_Z_R 0.1

module MUX81HSP (Z, D0, D1, D2, D3, D4, D5, D6, D7, A, B, C);

   output Z;
   input D0;
   input D1;
   input D2;
   input D3;
   input D4;
   input D5;
   input D6;
   input D7;
   input A;
   input B;
   input C;


   // gate-level netlist replaced by UDPs - 19 DEC 1995
   U_MUX4    u0 (OUT_UDP_D0_TO_3_IN, D0, D1, D2, D3, A, B);
   U_MUX4    u1 (OUT_UDP_D4_TO_7_IN, D4, D5, D6, D7, A, B);
   U_MUX2  u2 (Z, OUT_UDP_D0_TO_3_IN, OUT_UDP_D4_TO_7_IN, C);

   buf u3 (D7T, D7);
   buf u4 (D6T, D6);
   buf u5 (D5T, D5);
   buf u6 (D4T, D4);
   buf u7 (D3T, D3);
   buf u8 (D2T, D2);
   buf u9 (D1T, D1);
   buf u10 (D0T, D0);
   buf u11 (CT, C);
   buf u12 (BT, B);
   buf u13 (AT, A);
 
`ifdef tristatecheck
always @(D0T or D1T or D2T or D3T or D4T or D5T or D6T or D7T or AT or BT or CT)
begin
case ({C,B,A})
3'b000 : if (D0 === 1'bz)
                $display ("WARNING: Cell MUX81HSP used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D0 = %b at time %d", A, B, C, D0, $time);
3'b001 : if (D1 === 1'bz)
                $display ("WARNING: Cell MUX81HSP used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D1 = %b at time %d", A, B, C, D1, $time);
3'b010 : if (D2 === 1'bz)
                $display ("WARNING: Cell MUX81HSP used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D2 = %b at time %d", A, B, C, D2, $time);
3'b011 : if (D3 === 1'bz)
                $display ("WARNING: Cell MUX81HSP used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D3 = %b at time %d", A, B, C, D3, $time);
3'b100 : if (D4 === 1'bz)
                $display ("WARNING: Cell MUX81HSP used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D4 = %b at time %d", A, B, C, D4, $time);
3'b101 : if (D5 === 1'bz)
                $display ("WARNING: Cell MUX81HSP used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D5 = %b at time %d", A, B, C, D5, $time);
3'b110 : if (D6 === 1'bz)
                $display ("WARNING: Cell MUX81HSP used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D6 = %b at time %d", A, B, C, D6, $time);
3'b111 : if (D7 === 1'bz)
                $display ("WARNING: Cell MUX81HSP used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D7 = %b at time %d", A, B, C, D7, $time);
default:;
endcase
if (((A === 1'bx) || (B === 1'bx) || (C === 1'bx)) && 
    ((D0 === 1'bz) || (D1 === 1'bz) || (D2 === 1'bz) || (D3 === 1'bz) || (D4 === 1'bz) || (D5 === 1'bz) || (D6 === 1'bz) || (D7 === 1'bz)))
begin
        $display ("WARNING: Cell MUX81HSP used in IDDQ unsafe mode at time %d", $time);
        $display ("         with inputs at A = %b, B = %b, C = %b, D0 = %b, D1 = %b, D2 = %b, D3 = %b, D4 = %b, D5 = %b, D6 = %b, D7 = %b", 
           A, B, C, D0, D1, D2, D3, D4, D5, D6, D7);
end
end
`endif


`ifdef functional
`else
   specify

      if (!D3 && D7 && A && B || !D2 && D6 && !A && B || !D1 && D5 && A && !B || !D0 && D4 && !A && !B) (C +=> Z) = (`MUX81HSP_C_R_Z_R,`MUX81HSP_C_F_Z_F);
      if (D3 && !D7 && A && B || D2 && !D6 && !A && B || D1 && !D5 && A && !B || D0 && !D4 && !A && !B) (C -=> Z) = (`MUX81HSP_C_F_Z_R,`MUX81HSP_C_R_Z_F);
      if (!D5 && D7 && A && C || !D4 && D6 && !A && C || !D1 && D3 && A && !C || !D0 && D2 && !A && !C) (B +=> Z) = (`MUX81HSP_B_R_Z_R,`MUX81HSP_B_F_Z_F);
      if (D5 && !D7 && A && C || D4 && !D6 && !A && C || D1 && !D3 && A && !C || D0 && !D2 && !A && !C) (B -=> Z) = (`MUX81HSP_B_F_Z_R,`MUX81HSP_B_R_Z_F);
      if (!D6 && D7 && B && C || !D4 && D5 && !B && C || !D2 && D3 && B && !C || !D0 && D1 && !B && !C) (A +=> Z) = (`MUX81HSP_A_R_Z_R,`MUX81HSP_A_F_Z_F);
      if (D6 && !D7 && B && C || D4 && !D5 && !B && C || D2 && !D3 && B && !C || D0 && !D1 && !B && !C) (A -=> Z) = (`MUX81HSP_A_F_Z_R,`MUX81HSP_A_R_Z_F);
      (D7 +=> Z) = (`MUX81HSP_D7_R_Z_R,`MUX81HSP_D7_F_Z_F);
      (D6 +=> Z) = (`MUX81HSP_D6_R_Z_R,`MUX81HSP_D6_F_Z_F);
      (D5 +=> Z) = (`MUX81HSP_D5_R_Z_R,`MUX81HSP_D5_F_Z_F);
      (D4 +=> Z) = (`MUX81HSP_D4_R_Z_R,`MUX81HSP_D4_F_Z_F);
      (D3 +=> Z) = (`MUX81HSP_D3_R_Z_R,`MUX81HSP_D3_F_Z_F);
      (D2 +=> Z) = (`MUX81HSP_D2_R_Z_R,`MUX81HSP_D2_F_Z_F);
      (D1 +=> Z) = (`MUX81HSP_D1_R_Z_R,`MUX81HSP_D1_F_Z_F);
      (D0 +=> Z) = (`MUX81HSP_D0_R_Z_R,`MUX81HSP_D0_F_Z_F);

   endspecify
`endif


endmodule // MUX81HSP

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
  
//  END
// Created from CVS on Date :1998/07/07 13:19:11 and Version :1.1 //
 
//  START
// CELL MUX81HSX4 

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define MUX81HSX4_C_F_Z_F 0.1
`define MUX81HSX4_C_R_Z_R 0.1
`define MUX81HSX4_C_F_Z_R 0.1
`define MUX81HSX4_C_R_Z_F 0.1
`define MUX81HSX4_B_F_Z_F 0.1
`define MUX81HSX4_B_R_Z_R 0.1
`define MUX81HSX4_B_F_Z_R 0.1
`define MUX81HSX4_B_R_Z_F 0.1
`define MUX81HSX4_A_F_Z_F 0.1
`define MUX81HSX4_A_R_Z_R 0.1
`define MUX81HSX4_A_F_Z_R 0.1
`define MUX81HSX4_A_R_Z_F 0.1
`define MUX81HSX4_D7_F_Z_F 0.1
`define MUX81HSX4_D7_R_Z_R 0.1
`define MUX81HSX4_D6_F_Z_F 0.1
`define MUX81HSX4_D6_R_Z_R 0.1
`define MUX81HSX4_D5_F_Z_F 0.1
`define MUX81HSX4_D5_R_Z_R 0.1
`define MUX81HSX4_D4_F_Z_F 0.1
`define MUX81HSX4_D4_R_Z_R 0.1
`define MUX81HSX4_D3_F_Z_F 0.1
`define MUX81HSX4_D3_R_Z_R 0.1
`define MUX81HSX4_D2_F_Z_F 0.1
`define MUX81HSX4_D2_R_Z_R 0.1
`define MUX81HSX4_D1_F_Z_F 0.1
`define MUX81HSX4_D1_R_Z_R 0.1
`define MUX81HSX4_D0_F_Z_F 0.1
`define MUX81HSX4_D0_R_Z_R 0.1

module MUX81HSX4 (Z, D0, D1, D2, D3, D4, D5, D6, D7, A, B, C);

   output Z;
   input D0;
   input D1;
   input D2;
   input D3;
   input D4;
   input D5;
   input D6;
   input D7;
   input A;
   input B;
   input C;


   // gate-level netlist replaced by UDPs - 19 DEC 1995
   U_MUX4    u0 (OUT_UDP_D0_TO_3_IN, D0, D1, D2, D3, A, B);
   U_MUX4    u1 (OUT_UDP_D4_TO_7_IN, D4, D5, D6, D7, A, B);
   U_MUX2  u2 (Z, OUT_UDP_D0_TO_3_IN, OUT_UDP_D4_TO_7_IN, C);

   buf u3 (D7T, D7);
   buf u4 (D6T, D6);
   buf u5 (D5T, D5);
   buf u6 (D4T, D4);
   buf u7 (D3T, D3);
   buf u8 (D2T, D2);
   buf u9 (D1T, D1);
   buf u10 (D0T, D0);
   buf u11 (CT, C);
   buf u12 (BT, B);
   buf u13 (AT, A);
 
`ifdef tristatecheck
always @(D0T or D1T or D2T or D3T or D4T or D5T or D6T or D7T or AT or BT or CT)
begin
case ({C,B,A})
3'b000 : if (D0 === 1'bz)
                $display ("WARNING: Cell MUX81HSX4 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D0 = %b at time %d", A, B, C, D0, $time);
3'b001 : if (D1 === 1'bz)
                $display ("WARNING: Cell MUX81HSX4 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D1 = %b at time %d", A, B, C, D1, $time);
3'b010 : if (D2 === 1'bz)
                $display ("WARNING: Cell MUX81HSX4 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D2 = %b at time %d", A, B, C, D2, $time);
3'b011 : if (D3 === 1'bz)
                $display ("WARNING: Cell MUX81HSX4 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D3 = %b at time %d", A, B, C, D3, $time);
3'b100 : if (D4 === 1'bz)
                $display ("WARNING: Cell MUX81HSX4 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D4 = %b at time %d", A, B, C, D4, $time);
3'b101 : if (D5 === 1'bz)
                $display ("WARNING: Cell MUX81HSX4 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D5 = %b at time %d", A, B, C, D5, $time);
3'b110 : if (D6 === 1'bz)
                $display ("WARNING: Cell MUX81HSX4 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D6 = %b at time %d", A, B, C, D6, $time);
3'b111 : if (D7 === 1'bz)
                $display ("WARNING: Cell MUX81HSX4 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D7 = %b at time %d", A, B, C, D7, $time);
default:;
endcase
if (((A === 1'bx) || (B === 1'bx) || (C === 1'bx)) && 
    ((D0 === 1'bz) || (D1 === 1'bz) || (D2 === 1'bz) || (D3 === 1'bz) || (D4 === 1'bz) || (D5 === 1'bz) || (D6 === 1'bz) || (D7 === 1'bz)))
begin
        $display ("WARNING: Cell MUX81HSX4 used in IDDQ unsafe mode at time %d", $time);
        $display ("         with inputs at A = %b, B = %b, C = %b, D0 = %b, D1 = %b, D2 = %b, D3 = %b, D4 = %b, D5 = %b, D6 = %b, D7 = %b", 
           A, B, C, D0, D1, D2, D3, D4, D5, D6, D7);
end
end
`endif


`ifdef functional
`else
   specify

      if (!D3 && D7 && A && B || !D2 && D6 && !A && B || !D1 && D5 && A && !B || !D0 && D4 && !A && !B) (C +=> Z) = (`MUX81HSX4_C_R_Z_R,`MUX81HSX4_C_F_Z_F);
      if (D3 && !D7 && A && B || D2 && !D6 && !A && B || D1 && !D5 && A && !B || D0 && !D4 && !A && !B) (C -=> Z) = (`MUX81HSX4_C_F_Z_R,`MUX81HSX4_C_R_Z_F);
      if (!D5 && D7 && A && C || !D4 && D6 && !A && C || !D1 && D3 && A && !C || !D0 && D2 && !A && !C) (B +=> Z) = (`MUX81HSX4_B_R_Z_R,`MUX81HSX4_B_F_Z_F);
      if (D5 && !D7 && A && C || D4 && !D6 && !A && C || D1 && !D3 && A && !C || D0 && !D2 && !A && !C) (B -=> Z) = (`MUX81HSX4_B_F_Z_R,`MUX81HSX4_B_R_Z_F);
      if (!D6 && D7 && B && C || !D4 && D5 && !B && C || !D2 && D3 && B && !C || !D0 && D1 && !B && !C) (A +=> Z) = (`MUX81HSX4_A_R_Z_R,`MUX81HSX4_A_F_Z_F);
      if (D6 && !D7 && B && C || D4 && !D5 && !B && C || D2 && !D3 && B && !C || D0 && !D1 && !B && !C) (A -=> Z) = (`MUX81HSX4_A_F_Z_R,`MUX81HSX4_A_R_Z_F);
      (D7 +=> Z) = (`MUX81HSX4_D7_R_Z_R,`MUX81HSX4_D7_F_Z_F);
      (D6 +=> Z) = (`MUX81HSX4_D6_R_Z_R,`MUX81HSX4_D6_F_Z_F);
      (D5 +=> Z) = (`MUX81HSX4_D5_R_Z_R,`MUX81HSX4_D5_F_Z_F);
      (D4 +=> Z) = (`MUX81HSX4_D4_R_Z_R,`MUX81HSX4_D4_F_Z_F);
      (D3 +=> Z) = (`MUX81HSX4_D3_R_Z_R,`MUX81HSX4_D3_F_Z_F);
      (D2 +=> Z) = (`MUX81HSX4_D2_R_Z_R,`MUX81HSX4_D2_F_Z_F);
      (D1 +=> Z) = (`MUX81HSX4_D1_R_Z_R,`MUX81HSX4_D1_F_Z_F);
      (D0 +=> Z) = (`MUX81HSX4_D0_R_Z_R,`MUX81HSX4_D0_F_Z_F);

   endspecify
`endif


endmodule // MUX81HSX4

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
  
//  END
// Created from CVS on Date :1998/07/07 13:19:11 and Version :1.1 //
 
//  START
// CELL MUX81NHS 

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define MUX81NHS_C_F_Z_F 0.1
`define MUX81NHS_C_R_Z_R 0.1
`define MUX81NHS_C_F_Z_R 0.1
`define MUX81NHS_C_R_Z_F 0.1
`define MUX81NHS_B_F_Z_F 0.1
`define MUX81NHS_B_R_Z_R 0.1
`define MUX81NHS_B_F_Z_R 0.1
`define MUX81NHS_B_R_Z_F 0.1
`define MUX81NHS_A_F_Z_F 0.1
`define MUX81NHS_A_R_Z_R 0.1
`define MUX81NHS_A_F_Z_R 0.1
`define MUX81NHS_A_R_Z_F 0.1
`define MUX81NHS_D7_F_Z_R 0.1
`define MUX81NHS_D7_R_Z_F 0.1
`define MUX81NHS_D6_F_Z_R 0.1
`define MUX81NHS_D6_R_Z_F 0.1
`define MUX81NHS_D5_F_Z_R 0.1
`define MUX81NHS_D5_R_Z_F 0.1
`define MUX81NHS_D4_F_Z_R 0.1
`define MUX81NHS_D4_R_Z_F 0.1
`define MUX81NHS_D3_F_Z_R 0.1
`define MUX81NHS_D3_R_Z_F 0.1
`define MUX81NHS_D2_F_Z_R 0.1
`define MUX81NHS_D2_R_Z_F 0.1
`define MUX81NHS_D1_F_Z_R 0.1
`define MUX81NHS_D1_R_Z_F 0.1
`define MUX81NHS_D0_F_Z_R 0.1
`define MUX81NHS_D0_R_Z_F 0.1

module MUX81NHS (Z, D0, D1, D2, D3, D4, D5, D6, D7, A, B, C);

   output Z;
   input D0;
   input D1;
   input D2;
   input D3;
   input D4;
   input D5;
   input D6;
   input D7;
   input A;
   input B;
   input C;


   // gate-level netlist replaced by UDPs - 19 DEC 1995
   U_MUX4    u0 (OUT_UDP_D0_TO_3_IN, D0, D1, D2, D3, A, B);
   U_MUX4    u1 (OUT_UDP_D4_TO_7_IN, D4, D5, D6, D7, A, B);
   U_MUX2  u2 (ZX, OUT_UDP_D0_TO_3_IN, OUT_UDP_D4_TO_7_IN, C);
   not  u14 (Z, ZX);

   buf u3 (D7T, D7);
   buf u4 (D6T, D6);
   buf u5 (D5T, D5);
   buf u6 (D4T, D4);
   buf u7 (D3T, D3);
   buf u8 (D2T, D2);
   buf u9 (D1T, D1);
   buf u10 (D0T, D0);
   buf u11 (CT, C);
   buf u12 (BT, B);
   buf u13 (AT, A);
 
`ifdef tristatecheck
always @(D0T or D1T or D2T or D3T or D4T or D5T or D6T or D7T or AT or BT or CT)
begin
case ({C,B,A})
3'b000 : if (D0 === 1'bz)
                $display ("WARNING: Cell MUX81NHS used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D0 = %b at time %d", A, B, C, D0, $time);
3'b001 : if (D1 === 1'bz)
                $display ("WARNING: Cell MUX81NHS used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D1 = %b at time %d", A, B, C, D1, $time);
3'b010 : if (D2 === 1'bz)
                $display ("WARNING: Cell MUX81NHS used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D2 = %b at time %d", A, B, C, D2, $time);
3'b011 : if (D3 === 1'bz)
                $display ("WARNING: Cell MUX81NHS used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D3 = %b at time %d", A, B, C, D3, $time);
3'b100 : if (D4 === 1'bz)
                $display ("WARNING: Cell MUX81NHS used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D4 = %b at time %d", A, B, C, D4, $time);
3'b101 : if (D5 === 1'bz)
                $display ("WARNING: Cell MUX81NHS used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D5 = %b at time %d", A, B, C, D5, $time);
3'b110 : if (D6 === 1'bz)
                $display ("WARNING: Cell MUX81NHS used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D6 = %b at time %d", A, B, C, D6, $time);
3'b111 : if (D7 === 1'bz)
                $display ("WARNING: Cell MUX81NHS used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D7 = %b at time %d", A, B, C, D7, $time);
default:;
endcase
if (((A === 1'bx) || (B === 1'bx) || (C === 1'bx)) && 
    ((D0 === 1'bz) || (D1 === 1'bz) || (D2 === 1'bz) || (D3 === 1'bz) || (D4 === 1'bz) || (D5 === 1'bz) || (D6 === 1'bz) || (D7 === 1'bz)))
begin
        $display ("WARNING: Cell MUX81NHS used in IDDQ unsafe mode at time %d", $time);
        $display ("         with inputs at A = %b, B = %b, C = %b, D0 = %b, D1 = %b, D2 = %b, D3 = %b, D4 = %b, D5 = %b, D6 = %b, D7 = %b", 
           A, B, C, D0, D1, D2, D3, D4, D5, D6, D7);
end
end
`endif


`ifdef functional
`else
   specify

      if (!D3 && D7 && A && B || !D2 && D6 && !A && B || !D1 && D5 && A && !B || !D0 && D4 && !A && !B) (C -=> Z) = (`MUX81NHS_C_F_Z_R,`MUX81NHS_C_R_Z_F);
      if (D3 && !D7 && A && B || D2 && !D6 && !A && B || D1 && !D5 && A && !B || D0 && !D4 && !A && !B) (C +=> Z) = (`MUX81NHS_C_R_Z_R,`MUX81NHS_C_F_Z_F);
      if (!D5 && D7 && A && C || !D4 && D6 && !A && C || !D1 && D3 && A && !C || !D0 && D2 && !A && !C) (B -=> Z) = (`MUX81NHS_B_F_Z_R,`MUX81NHS_B_R_Z_F);
      if (D5 && !D7 && A && C || D4 && !D6 && !A && C || D1 && !D3 && A && !C || D0 && !D2 && !A && !C) (B +=> Z) = (`MUX81NHS_B_R_Z_R,`MUX81NHS_B_F_Z_F);
      if (!D6 && D7 && B && C || !D4 && D5 && !B && C || !D2 && D3 && B && !C || !D0 && D1 && !B && !C) (A -=> Z) = (`MUX81NHS_A_F_Z_R,`MUX81NHS_A_R_Z_F);
      if (D6 && !D7 && B && C || D4 && !D5 && !B && C || D2 && !D3 && B && !C || D0 && !D1 && !B && !C) (A +=> Z) = (`MUX81NHS_A_R_Z_R,`MUX81NHS_A_F_Z_F);
      (D7 -=> Z) = (`MUX81NHS_D7_F_Z_R,`MUX81NHS_D7_R_Z_F);
      (D6 -=> Z) = (`MUX81NHS_D6_F_Z_R,`MUX81NHS_D6_R_Z_F);
      (D5 -=> Z) = (`MUX81NHS_D5_F_Z_R,`MUX81NHS_D5_R_Z_F);
      (D4 -=> Z) = (`MUX81NHS_D4_F_Z_R,`MUX81NHS_D4_R_Z_F);
      (D3 -=> Z) = (`MUX81NHS_D3_F_Z_R,`MUX81NHS_D3_R_Z_F);
      (D2 -=> Z) = (`MUX81NHS_D2_F_Z_R,`MUX81NHS_D2_R_Z_F);
      (D1 -=> Z) = (`MUX81NHS_D1_F_Z_R,`MUX81NHS_D1_R_Z_F);
      (D0 -=> Z) = (`MUX81NHS_D0_F_Z_R,`MUX81NHS_D0_R_Z_F);

   endspecify
`endif


endmodule // MUX81NHS

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
//  END
// Created from CVS on Date :1998/07/07 13:19:11 and Version :1.1 //
 
//  START
// CELL MUX81NHSP 

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define MUX81NHSP_C_F_Z_F 0.1
`define MUX81NHSP_C_R_Z_R 0.1
`define MUX81NHSP_C_F_Z_R 0.1
`define MUX81NHSP_C_R_Z_F 0.1
`define MUX81NHSP_B_F_Z_F 0.1
`define MUX81NHSP_B_R_Z_R 0.1
`define MUX81NHSP_B_F_Z_R 0.1
`define MUX81NHSP_B_R_Z_F 0.1
`define MUX81NHSP_A_F_Z_F 0.1
`define MUX81NHSP_A_R_Z_R 0.1
`define MUX81NHSP_A_F_Z_R 0.1
`define MUX81NHSP_A_R_Z_F 0.1
`define MUX81NHSP_D7_F_Z_R 0.1
`define MUX81NHSP_D7_R_Z_F 0.1
`define MUX81NHSP_D6_F_Z_R 0.1
`define MUX81NHSP_D6_R_Z_F 0.1
`define MUX81NHSP_D5_F_Z_R 0.1
`define MUX81NHSP_D5_R_Z_F 0.1
`define MUX81NHSP_D4_F_Z_R 0.1
`define MUX81NHSP_D4_R_Z_F 0.1
`define MUX81NHSP_D3_F_Z_R 0.1
`define MUX81NHSP_D3_R_Z_F 0.1
`define MUX81NHSP_D2_F_Z_R 0.1
`define MUX81NHSP_D2_R_Z_F 0.1
`define MUX81NHSP_D1_F_Z_R 0.1
`define MUX81NHSP_D1_R_Z_F 0.1
`define MUX81NHSP_D0_F_Z_R 0.1
`define MUX81NHSP_D0_R_Z_F 0.1

module MUX81NHSP (Z, D0, D1, D2, D3, D4, D5, D6, D7, A, B, C);

   output Z;
   input D0;
   input D1;
   input D2;
   input D3;
   input D4;
   input D5;
   input D6;
   input D7;
   input A;
   input B;
   input C;


   // gate-level netlist replaced by UDPs - 19 DEC 1995
   U_MUX4    u0 (OUT_UDP_D0_TO_3_IN, D0, D1, D2, D3, A, B);
   U_MUX4    u1 (OUT_UDP_D4_TO_7_IN, D4, D5, D6, D7, A, B);
   U_MUX2  u2 (ZX, OUT_UDP_D0_TO_3_IN, OUT_UDP_D4_TO_7_IN, C);
   not  u14 (Z, ZX);

   buf u3 (D7T, D7);
   buf u4 (D6T, D6);
   buf u5 (D5T, D5);
   buf u6 (D4T, D4);
   buf u7 (D3T, D3);
   buf u8 (D2T, D2);
   buf u9 (D1T, D1);
   buf u10 (D0T, D0);
   buf u11 (CT, C);
   buf u12 (BT, B);
   buf u13 (AT, A);
 
`ifdef tristatecheck
always @(D0T or D1T or D2T or D3T or D4T or D5T or D6T or D7T or AT or BT or CT)
begin
case ({C,B,A})
3'b000 : if (D0 === 1'bz)
                $display ("WARNING: Cell MUX81NHSP used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D0 = %b at time %d", A, B, C, D0, $time);
3'b001 : if (D1 === 1'bz)
                $display ("WARNING: Cell MUX81NHSP used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D1 = %b at time %d", A, B, C, D1, $time);
3'b010 : if (D2 === 1'bz)
                $display ("WARNING: Cell MUX81NHSP used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D2 = %b at time %d", A, B, C, D2, $time);
3'b011 : if (D3 === 1'bz)
                $display ("WARNING: Cell MUX81NHSP used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D3 = %b at time %d", A, B, C, D3, $time);
3'b100 : if (D4 === 1'bz)
                $display ("WARNING: Cell MUX81NHSP used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D4 = %b at time %d", A, B, C, D4, $time);
3'b101 : if (D5 === 1'bz)
                $display ("WARNING: Cell MUX81NHSP used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D5 = %b at time %d", A, B, C, D5, $time);
3'b110 : if (D6 === 1'bz)
                $display ("WARNING: Cell MUX81NHSP used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D6 = %b at time %d", A, B, C, D6, $time);
3'b111 : if (D7 === 1'bz)
                $display ("WARNING: Cell MUX81NHSP used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D7 = %b at time %d", A, B, C, D7, $time);
default:;
endcase
if (((A === 1'bx) || (B === 1'bx) || (C === 1'bx)) && 
    ((D0 === 1'bz) || (D1 === 1'bz) || (D2 === 1'bz) || (D3 === 1'bz) || (D4 === 1'bz) || (D5 === 1'bz) || (D6 === 1'bz) || (D7 === 1'bz)))
begin
        $display ("WARNING: Cell MUX81NHSP used in IDDQ unsafe mode at time %d", $time);
        $display ("         with inputs at A = %b, B = %b, C = %b, D0 = %b, D1 = %b, D2 = %b, D3 = %b, D4 = %b, D5 = %b, D6 = %b, D7 = %b", 
           A, B, C, D0, D1, D2, D3, D4, D5, D6, D7);
end
end
`endif


`ifdef functional
`else
   specify

      if (!D3 && D7 && A && B || !D2 && D6 && !A && B || !D1 && D5 && A && !B || !D0 && D4 && !A && !B) (C -=> Z) = (`MUX81NHSP_C_F_Z_R,`MUX81NHSP_C_R_Z_F);
      if (D3 && !D7 && A && B || D2 && !D6 && !A && B || D1 && !D5 && A && !B || D0 && !D4 && !A && !B) (C +=> Z) = (`MUX81NHSP_C_R_Z_R,`MUX81NHSP_C_F_Z_F);
      if (!D5 && D7 && A && C || !D4 && D6 && !A && C || !D1 && D3 && A && !C || !D0 && D2 && !A && !C) (B -=> Z) = (`MUX81NHSP_B_F_Z_R,`MUX81NHSP_B_R_Z_F);
      if (D5 && !D7 && A && C || D4 && !D6 && !A && C || D1 && !D3 && A && !C || D0 && !D2 && !A && !C) (B +=> Z) = (`MUX81NHSP_B_R_Z_R,`MUX81NHSP_B_F_Z_F);
      if (!D6 && D7 && B && C || !D4 && D5 && !B && C || !D2 && D3 && B && !C || !D0 && D1 && !B && !C) (A -=> Z) = (`MUX81NHSP_A_F_Z_R,`MUX81NHSP_A_R_Z_F);
      if (D6 && !D7 && B && C || D4 && !D5 && !B && C || D2 && !D3 && B && !C || D0 && !D1 && !B && !C) (A +=> Z) = (`MUX81NHSP_A_R_Z_R,`MUX81NHSP_A_F_Z_F);
      (D7 -=> Z) = (`MUX81NHSP_D7_F_Z_R,`MUX81NHSP_D7_R_Z_F);
      (D6 -=> Z) = (`MUX81NHSP_D6_F_Z_R,`MUX81NHSP_D6_R_Z_F);
      (D5 -=> Z) = (`MUX81NHSP_D5_F_Z_R,`MUX81NHSP_D5_R_Z_F);
      (D4 -=> Z) = (`MUX81NHSP_D4_F_Z_R,`MUX81NHSP_D4_R_Z_F);
      (D3 -=> Z) = (`MUX81NHSP_D3_F_Z_R,`MUX81NHSP_D3_R_Z_F);
      (D2 -=> Z) = (`MUX81NHSP_D2_F_Z_R,`MUX81NHSP_D2_R_Z_F);
      (D1 -=> Z) = (`MUX81NHSP_D1_F_Z_R,`MUX81NHSP_D1_R_Z_F);
      (D0 -=> Z) = (`MUX81NHSP_D0_F_Z_R,`MUX81NHSP_D0_R_Z_F);

   endspecify
`endif


endmodule // MUX81NHSP

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
//  END
// Created from CVS on Date :1998/07/07 13:19:11 and Version :1.1 //
 
//  START
// CELL MUX81NHSX4 

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif

`define MUX81NHSX4_C_F_Z_F 0.1
`define MUX81NHSX4_C_R_Z_R 0.1
`define MUX81NHSX4_C_F_Z_R 0.1
`define MUX81NHSX4_C_R_Z_F 0.1
`define MUX81NHSX4_B_F_Z_F 0.1
`define MUX81NHSX4_B_R_Z_R 0.1
`define MUX81NHSX4_B_F_Z_R 0.1
`define MUX81NHSX4_B_R_Z_F 0.1
`define MUX81NHSX4_A_F_Z_F 0.1
`define MUX81NHSX4_A_R_Z_R 0.1
`define MUX81NHSX4_A_F_Z_R 0.1
`define MUX81NHSX4_A_R_Z_F 0.1
`define MUX81NHSX4_D7_F_Z_R 0.1
`define MUX81NHSX4_D7_R_Z_F 0.1
`define MUX81NHSX4_D6_F_Z_R 0.1
`define MUX81NHSX4_D6_R_Z_F 0.1
`define MUX81NHSX4_D5_F_Z_R 0.1
`define MUX81NHSX4_D5_R_Z_F 0.1
`define MUX81NHSX4_D4_F_Z_R 0.1
`define MUX81NHSX4_D4_R_Z_F 0.1
`define MUX81NHSX4_D3_F_Z_R 0.1
`define MUX81NHSX4_D3_R_Z_F 0.1
`define MUX81NHSX4_D2_F_Z_R 0.1
`define MUX81NHSX4_D2_R_Z_F 0.1
`define MUX81NHSX4_D1_F_Z_R 0.1
`define MUX81NHSX4_D1_R_Z_F 0.1
`define MUX81NHSX4_D0_F_Z_R 0.1
`define MUX81NHSX4_D0_R_Z_F 0.1

module MUX81NHSX4 (Z, D0, D1, D2, D3, D4, D5, D6, D7, A, B, C);

   output Z;
   input D0;
   input D1;
   input D2;
   input D3;
   input D4;
   input D5;
   input D6;
   input D7;
   input A;
   input B;
   input C;


   // gate-level netlist replaced by UDPs - 19 DEC 1995
   U_MUX4    u0 (OUT_UDP_D0_TO_3_IN, D0, D1, D2, D3, A, B);
   U_MUX4    u1 (OUT_UDP_D4_TO_7_IN, D4, D5, D6, D7, A, B);
   U_MUX2  u2 (ZX, OUT_UDP_D0_TO_3_IN, OUT_UDP_D4_TO_7_IN, C);
   not  u14 (Z, ZX);

   buf u3 (D7T, D7);
   buf u4 (D6T, D6);
   buf u5 (D5T, D5);
   buf u6 (D4T, D4);
   buf u7 (D3T, D3);
   buf u8 (D2T, D2);
   buf u9 (D1T, D1);
   buf u10 (D0T, D0);
   buf u11 (CT, C);
   buf u12 (BT, B);
   buf u13 (AT, A);
 
`ifdef tristatecheck
always @(D0T or D1T or D2T or D3T or D4T or D5T or D6T or D7T or AT or BT or CT)
begin
case ({C,B,A})
3'b000 : if (D0 === 1'bz)
                $display ("WARNING: Cell MUX81NHSX4 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D0 = %b at time %d", A, B, C, D0, $time);
3'b001 : if (D1 === 1'bz)
                $display ("WARNING: Cell MUX81NHSX4 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D1 = %b at time %d", A, B, C, D1, $time);
3'b010 : if (D2 === 1'bz)
                $display ("WARNING: Cell MUX81NHSX4 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D2 = %b at time %d", A, B, C, D2, $time);
3'b011 : if (D3 === 1'bz)
                $display ("WARNING: Cell MUX81NHSX4 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D3 = %b at time %d", A, B, C, D3, $time);
3'b100 : if (D4 === 1'bz)
                $display ("WARNING: Cell MUX81NHSX4 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D4 = %b at time %d", A, B, C, D4, $time);
3'b101 : if (D5 === 1'bz)
                $display ("WARNING: Cell MUX81NHSX4 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D5 = %b at time %d", A, B, C, D5, $time);
3'b110 : if (D6 === 1'bz)
                $display ("WARNING: Cell MUX81NHSX4 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D6 = %b at time %d", A, B, C, D6, $time);
3'b111 : if (D7 === 1'bz)
                $display ("WARNING: Cell MUX81NHSX4 used in IDDQ unsafe mode with A = %b, B = %b, C = %b, D7 = %b at time %d", A, B, C, D7, $time);
default:;
endcase
if (((A === 1'bx) || (B === 1'bx) || (C === 1'bx)) && 
    ((D0 === 1'bz) || (D1 === 1'bz) || (D2 === 1'bz) || (D3 === 1'bz) || (D4 === 1'bz) || (D5 === 1'bz) || (D6 === 1'bz) || (D7 === 1'bz)))
begin
        $display ("WARNING: Cell MUX81NHSX4 used in IDDQ unsafe mode at time %d", $time);
        $display ("         with inputs at A = %b, B = %b, C = %b, D0 = %b, D1 = %b, D2 = %b, D3 = %b, D4 = %b, D5 = %b, D6 = %b, D7 = %b", 
           A, B, C, D0, D1, D2, D3, D4, D5, D6, D7);
end
end
`endif


`ifdef functional
`else
   specify

      if (!D3 && D7 && A && B || !D2 && D6 && !A && B || !D1 && D5 && A && !B || !D0 && D4 && !A && !B) (C -=> Z) = (`MUX81NHSX4_C_F_Z_R,`MUX81NHSX4_C_R_Z_F);
      if (D3 && !D7 && A && B || D2 && !D6 && !A && B || D1 && !D5 && A && !B || D0 && !D4 && !A && !B) (C +=> Z) = (`MUX81NHSX4_C_R_Z_R,`MUX81NHSX4_C_F_Z_F);
      if (!D5 && D7 && A && C || !D4 && D6 && !A && C || !D1 && D3 && A && !C || !D0 && D2 && !A && !C) (B -=> Z) = (`MUX81NHSX4_B_F_Z_R,`MUX81NHSX4_B_R_Z_F);
      if (D5 && !D7 && A && C || D4 && !D6 && !A && C || D1 && !D3 && A && !C || D0 && !D2 && !A && !C) (B +=> Z) = (`MUX81NHSX4_B_R_Z_R,`MUX81NHSX4_B_F_Z_F);
      if (!D6 && D7 && B && C || !D4 && D5 && !B && C || !D2 && D3 && B && !C || !D0 && D1 && !B && !C) (A -=> Z) = (`MUX81NHSX4_A_F_Z_R,`MUX81NHSX4_A_R_Z_F);
      if (D6 && !D7 && B && C || D4 && !D5 && !B && C || D2 && !D3 && B && !C || D0 && !D1 && !B && !C) (A +=> Z) = (`MUX81NHSX4_A_R_Z_R,`MUX81NHSX4_A_F_Z_F);
      (D7 -=> Z) = (`MUX81NHSX4_D7_F_Z_R,`MUX81NHSX4_D7_R_Z_F);
      (D6 -=> Z) = (`MUX81NHSX4_D6_F_Z_R,`MUX81NHSX4_D6_R_Z_F);
      (D5 -=> Z) = (`MUX81NHSX4_D5_F_Z_R,`MUX81NHSX4_D5_R_Z_F);
      (D4 -=> Z) = (`MUX81NHSX4_D4_F_Z_R,`MUX81NHSX4_D4_R_Z_F);
      (D3 -=> Z) = (`MUX81NHSX4_D3_F_Z_R,`MUX81NHSX4_D3_R_Z_F);
      (D2 -=> Z) = (`MUX81NHSX4_D2_F_Z_R,`MUX81NHSX4_D2_R_Z_F);
      (D1 -=> Z) = (`MUX81NHSX4_D1_F_Z_R,`MUX81NHSX4_D1_R_Z_F);
      (D0 -=> Z) = (`MUX81NHSX4_D0_F_Z_R,`MUX81NHSX4_D0_R_Z_F);

   endspecify
`endif


endmodule // MUX81NHSX4

`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine
 
//  END
// Created from CVS on Date :1998/07/07 13:19:11 and Version :1.1 //
 
//  START
// CELL ND2HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND2HSX05_B_F_Z_R 0.1
`define ND2HSX05_B_R_Z_F 0.1
`define ND2HSX05_A_F_Z_R 0.1
`define ND2HSX05_A_R_Z_F 0.1

module ND2HSX05 (Z, A, B);

   output Z;
   input A;
   input B;


   nand  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`ND2HSX05_B_F_Z_R,`ND2HSX05_B_R_Z_F);
      (A -=> Z) = (`ND2HSX05_A_F_Z_R,`ND2HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // ND2HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:22 and Version :1.1 //
 
//  START 
// CELL ND2HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND2HS_B_F_Z_R 0.1
`define ND2HS_B_R_Z_F 0.1
`define ND2HS_A_F_Z_R 0.1
`define ND2HS_A_R_Z_F 0.1

module ND2HS (Z, A, B);

   output Z;
   input A;
   input B;


   nand  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`ND2HS_B_F_Z_R,`ND2HS_B_R_Z_F);
      (A -=> Z) = (`ND2HS_A_F_Z_R,`ND2HS_A_R_Z_F);

   endspecify
`endif


endmodule // ND2HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:22 and Version :1.1 //
 
//  START 
// CELL ND2HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND2HSP_B_F_Z_R 0.1
`define ND2HSP_B_R_Z_F 0.1
`define ND2HSP_A_F_Z_R 0.1
`define ND2HSP_A_R_Z_F 0.1

module ND2HSP (Z, A, B);

   output Z;
   input A;
   input B;


   nand  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`ND2HSP_B_F_Z_R,`ND2HSP_B_R_Z_F);
      (A -=> Z) = (`ND2HSP_A_F_Z_R,`ND2HSP_A_R_Z_F);

   endspecify
`endif


endmodule // ND2HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:22 and Version :1.1 //
 
//  START 
// CELL ND2HSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND2HSX3_B_F_Z_R 0.1
`define ND2HSX3_B_R_Z_F 0.1
`define ND2HSX3_A_F_Z_R 0.1
`define ND2HSX3_A_R_Z_F 0.1

module ND2HSX3 (Z, A, B);

   output Z;
   input A;
   input B;


   nand  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`ND2HSX3_B_F_Z_R,`ND2HSX3_B_R_Z_F);
      (A -=> Z) = (`ND2HSX3_A_F_Z_R,`ND2HSX3_A_R_Z_F);

   endspecify
`endif


endmodule // ND2HSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:22 and Version :1.1 //
 
//  START 
// CELL ND2HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND2HSX4_B_F_Z_R 0.1
`define ND2HSX4_B_R_Z_F 0.1
`define ND2HSX4_A_F_Z_R 0.1
`define ND2HSX4_A_R_Z_F 0.1

module ND2HSX4 (Z, A, B);

   output Z;
   input A;
   input B;


   nand  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`ND2HSX4_B_F_Z_R,`ND2HSX4_B_R_Z_F);
      (A -=> Z) = (`ND2HSX4_A_F_Z_R,`ND2HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // ND2HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:22 and Version :1.1 //
 
//  START 
// CELL B_ND2HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define B_ND2HSX4_B_F_Z_R 0.1
`define B_ND2HSX4_B_R_Z_F 0.1
`define B_ND2HSX4_A_F_Z_R 0.1
`define B_ND2HSX4_A_R_Z_F 0.1

module B_ND2HSX4 (Z, A, B);

   output Z;
   input A;
   input B;


   nand  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`B_ND2HSX4_B_F_Z_R,`B_ND2HSX4_B_R_Z_F);
      (A -=> Z) = (`B_ND2HSX4_A_F_Z_R,`B_ND2HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // B_ND2HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:22 and Version :1.1 //
 
//  START 
// CELL F_ND2HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_ND2HSX4_B_F_Z_R 0.1
`define F_ND2HSX4_B_R_Z_F 0.1
`define F_ND2HSX4_A_F_Z_R 0.1
`define F_ND2HSX4_A_R_Z_F 0.1

module F_ND2HSX4 (Z, A, B);

   output Z;
   input A;
   input B;


   nand  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`F_ND2HSX4_B_F_Z_R,`F_ND2HSX4_B_R_Z_F);
      (A -=> Z) = (`F_ND2HSX4_A_F_Z_R,`F_ND2HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // F_ND2HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:22 and Version :1.1 //
 
//  START 
// CELL F_ND2HSX6

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_ND2HSX6_B_F_Z_R 0.1
`define F_ND2HSX6_B_R_Z_F 0.1
`define F_ND2HSX6_A_F_Z_R 0.1
`define F_ND2HSX6_A_R_Z_F 0.1

module F_ND2HSX6 (Z, A, B);

   output Z;
   input A;
   input B;


   nand  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`F_ND2HSX6_B_F_Z_R,`F_ND2HSX6_B_R_Z_F);
      (A -=> Z) = (`F_ND2HSX6_A_F_Z_R,`F_ND2HSX6_A_R_Z_F);

   endspecify
`endif


endmodule // F_ND2HSX6
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:22 and Version :1.1 //
 
//  START 
// CELL F_ND2HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_ND2HSX8_B_F_Z_R 0.1
`define F_ND2HSX8_B_R_Z_F 0.1
`define F_ND2HSX8_A_F_Z_R 0.1
`define F_ND2HSX8_A_R_Z_F 0.1

module F_ND2HSX8 (Z, A, B);

   output Z;
   input A;
   input B;


   nand  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`F_ND2HSX8_B_F_Z_R,`F_ND2HSX8_B_R_Z_F);
      (A -=> Z) = (`F_ND2HSX8_A_F_Z_R,`F_ND2HSX8_A_R_Z_F);

   endspecify
`endif


endmodule // F_ND2HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:22 and Version :1.1 //
 
//  START 
// CELL M_ND2HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define M_ND2HSP_B_F_Z_R 0.1
`define M_ND2HSP_B_R_Z_F 0.1
`define M_ND2HSP_A_F_Z_R 0.1
`define M_ND2HSP_A_R_Z_F 0.1

module M_ND2HSP (Z, A, B);

   output Z;
   input A;
   input B;


   nand  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`M_ND2HSP_B_F_Z_R,`M_ND2HSP_B_R_Z_F);
      (A -=> Z) = (`M_ND2HSP_A_F_Z_R,`M_ND2HSP_A_R_Z_F);

   endspecify
`endif


endmodule // M_ND2HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:22 and Version :1.1 //
 
//  START 
// CELL M_ND2HSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define M_ND2HSX3_B_F_Z_R 0.1
`define M_ND2HSX3_B_R_Z_F 0.1
`define M_ND2HSX3_A_F_Z_R 0.1
`define M_ND2HSX3_A_R_Z_F 0.1

module M_ND2HSX3 (Z, A, B);

   output Z;
   input A;
   input B;


   nand  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`M_ND2HSX3_B_F_Z_R,`M_ND2HSX3_B_R_Z_F);
      (A -=> Z) = (`M_ND2HSX3_A_F_Z_R,`M_ND2HSX3_A_R_Z_F);

   endspecify
`endif


endmodule // M_ND2HSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:22 and Version :1.1 //
 
//  START 
// CELL ND2AHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND2AHS_B_F_Z_R 0.1
`define ND2AHS_B_R_Z_F 0.1
`define ND2AHS_A_F_Z_F 0.1
`define ND2AHS_A_R_Z_R 0.1

module ND2AHS (Z, A, B);

   output Z;
   input A;
   input B;


   or  u0 (Z, A, BX);
   not  u1 (BX, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`ND2AHS_B_F_Z_R,`ND2AHS_B_R_Z_F);
      (A +=> Z) = (`ND2AHS_A_R_Z_R,`ND2AHS_A_F_Z_F);

   endspecify
`endif


endmodule // ND2AHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:22 and Version :1.1 //
 
//  START 
// CELL ND2AHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND2AHSP_B_F_Z_R 0.1
`define ND2AHSP_B_R_Z_F 0.1
`define ND2AHSP_A_F_Z_F 0.1
`define ND2AHSP_A_R_Z_R 0.1

module ND2AHSP (Z, A, B);

   output Z;
   input A;
   input B;


   or  u0 (Z, A, BX);
   not  u1 (BX, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`ND2AHSP_B_F_Z_R,`ND2AHSP_B_R_Z_F);
      (A +=> Z) = (`ND2AHSP_A_R_Z_R,`ND2AHSP_A_F_Z_F);

   endspecify
`endif


endmodule // ND2AHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:22 and Version :1.1 //
 
//  START 
// CELL ND2AHSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND2AHSX3_B_F_Z_R 0.1
`define ND2AHSX3_B_R_Z_F 0.1
`define ND2AHSX3_A_F_Z_F 0.1
`define ND2AHSX3_A_R_Z_R 0.1

module ND2AHSX3 (Z, A, B);

   output Z;
   input A;
   input B;


   or  u0 (Z, A, BX);
   not  u1 (BX, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`ND2AHSX3_B_F_Z_R,`ND2AHSX3_B_R_Z_F);
      (A +=> Z) = (`ND2AHSX3_A_R_Z_R,`ND2AHSX3_A_F_Z_F);

   endspecify
`endif


endmodule // ND2AHSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:22 and Version :1.1 //
 
//  START 
// CELL ND2AHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND2AHSX4_B_F_Z_R 0.1
`define ND2AHSX4_B_R_Z_F 0.1
`define ND2AHSX4_A_F_Z_F 0.1
`define ND2AHSX4_A_R_Z_R 0.1

module ND2AHSX4 (Z, A, B);

   output Z;
   input A;
   input B;


   or  u0 (Z, A, BX);
   not  u1 (BX, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`ND2AHSX4_B_F_Z_R,`ND2AHSX4_B_R_Z_F);
      (A +=> Z) = (`ND2AHSX4_A_R_Z_R,`ND2AHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // ND2AHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:22 and Version :1.1 //
 
//  START 
// CELL F_ND2AHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_ND2AHSP_B_F_Z_R 0.1
`define F_ND2AHSP_B_R_Z_F 0.1
`define F_ND2AHSP_A_F_Z_F 0.1
`define F_ND2AHSP_A_R_Z_R 0.1

module F_ND2AHSP (Z, A, B);

   output Z;
   input A;
   input B;


   or  u0 (Z, A, BX);
   not  u1 (BX, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`F_ND2AHSP_B_F_Z_R,`F_ND2AHSP_B_R_Z_F);
      (A +=> Z) = (`F_ND2AHSP_A_R_Z_R,`F_ND2AHSP_A_F_Z_F);

   endspecify
`endif


endmodule // F_ND2AHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:22 and Version :1.1 //
 
//  START 
// CELL F_ND2AHSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_ND2AHSX3_B_F_Z_R 0.1
`define F_ND2AHSX3_B_R_Z_F 0.1
`define F_ND2AHSX3_A_F_Z_F 0.1
`define F_ND2AHSX3_A_R_Z_R 0.1

module F_ND2AHSX3 (Z, A, B);

   output Z;
   input A;
   input B;


   or  u0 (Z, A, BX);
   not  u1 (BX, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`F_ND2AHSX3_B_F_Z_R,`F_ND2AHSX3_B_R_Z_F);
      (A +=> Z) = (`F_ND2AHSX3_A_R_Z_R,`F_ND2AHSX3_A_F_Z_F);

   endspecify
`endif


endmodule // F_ND2AHSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:22 and Version :1.1 //
 
//  START 
// CELL F_ND2AHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_ND2AHSX4_B_F_Z_R 0.1
`define F_ND2AHSX4_B_R_Z_F 0.1
`define F_ND2AHSX4_A_F_Z_F 0.1
`define F_ND2AHSX4_A_R_Z_R 0.1

module F_ND2AHSX4 (Z, A, B);

   output Z;
   input A;
   input B;


   or  u0 (Z, A, BX);
   not  u1 (BX, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`F_ND2AHSX4_B_F_Z_R,`F_ND2AHSX4_B_R_Z_F);
      (A +=> Z) = (`F_ND2AHSX4_A_R_Z_R,`F_ND2AHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // F_ND2AHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:22 and Version :1.1 //
 
//  START 
// CELL F_ND2AHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_ND2AHSX8_B_F_Z_R 0.1
`define F_ND2AHSX8_B_R_Z_F 0.1
`define F_ND2AHSX8_A_F_Z_F 0.1
`define F_ND2AHSX8_A_R_Z_R 0.1

module F_ND2AHSX8 (Z, A, B);

   output Z;
   input A;
   input B;


   or  u0 (Z, A, BX);
   not  u1 (BX, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`F_ND2AHSX8_B_F_Z_R,`F_ND2AHSX8_B_R_Z_F);
      (A +=> Z) = (`F_ND2AHSX8_A_R_Z_R,`F_ND2AHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // F_ND2AHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:22 and Version :1.1 //
 
//  START 
// CELL ND3HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND3HSX05_C_F_Z_R 0.1
`define ND3HSX05_C_R_Z_F 0.1
`define ND3HSX05_B_F_Z_R 0.1
`define ND3HSX05_B_R_Z_F 0.1
`define ND3HSX05_A_F_Z_R 0.1
`define ND3HSX05_A_R_Z_F 0.1

module ND3HSX05 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C -=> Z) = (`ND3HSX05_C_F_Z_R,`ND3HSX05_C_R_Z_F);
      (B -=> Z) = (`ND3HSX05_B_F_Z_R,`ND3HSX05_B_R_Z_F);
      (A -=> Z) = (`ND3HSX05_A_F_Z_R,`ND3HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // ND3HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:29 and Version :1.1 //
 
//  START 
// CELL ND3HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND3HS_C_F_Z_R 0.1
`define ND3HS_C_R_Z_F 0.1
`define ND3HS_B_F_Z_R 0.1
`define ND3HS_B_R_Z_F 0.1
`define ND3HS_A_F_Z_R 0.1
`define ND3HS_A_R_Z_F 0.1

module ND3HS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C -=> Z) = (`ND3HS_C_F_Z_R,`ND3HS_C_R_Z_F);
      (B -=> Z) = (`ND3HS_B_F_Z_R,`ND3HS_B_R_Z_F);
      (A -=> Z) = (`ND3HS_A_F_Z_R,`ND3HS_A_R_Z_F);

   endspecify
`endif


endmodule // ND3HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:29 and Version :1.1 //
 
//  START 
// CELL ND3HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND3HSP_C_F_Z_R 0.1
`define ND3HSP_C_R_Z_F 0.1
`define ND3HSP_B_F_Z_R 0.1
`define ND3HSP_B_R_Z_F 0.1
`define ND3HSP_A_F_Z_R 0.1
`define ND3HSP_A_R_Z_F 0.1

module ND3HSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C -=> Z) = (`ND3HSP_C_F_Z_R,`ND3HSP_C_R_Z_F);
      (B -=> Z) = (`ND3HSP_B_F_Z_R,`ND3HSP_B_R_Z_F);
      (A -=> Z) = (`ND3HSP_A_F_Z_R,`ND3HSP_A_R_Z_F);

   endspecify
`endif


endmodule // ND3HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:29 and Version :1.1 //
 
//  START 
// CELL ND3HSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND3HSX3_C_F_Z_R 0.1
`define ND3HSX3_C_R_Z_F 0.1
`define ND3HSX3_B_F_Z_R 0.1
`define ND3HSX3_B_R_Z_F 0.1
`define ND3HSX3_A_F_Z_R 0.1
`define ND3HSX3_A_R_Z_F 0.1

module ND3HSX3 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C -=> Z) = (`ND3HSX3_C_F_Z_R,`ND3HSX3_C_R_Z_F);
      (B -=> Z) = (`ND3HSX3_B_F_Z_R,`ND3HSX3_B_R_Z_F);
      (A -=> Z) = (`ND3HSX3_A_F_Z_R,`ND3HSX3_A_R_Z_F);

   endspecify
`endif


endmodule // ND3HSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:29 and Version :1.1 //
 
//  START 
// CELL ND3HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND3HSX4_C_F_Z_R 0.1
`define ND3HSX4_C_R_Z_F 0.1
`define ND3HSX4_B_F_Z_R 0.1
`define ND3HSX4_B_R_Z_F 0.1
`define ND3HSX4_A_F_Z_R 0.1
`define ND3HSX4_A_R_Z_F 0.1

module ND3HSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C -=> Z) = (`ND3HSX4_C_F_Z_R,`ND3HSX4_C_R_Z_F);
      (B -=> Z) = (`ND3HSX4_B_F_Z_R,`ND3HSX4_B_R_Z_F);
      (A -=> Z) = (`ND3HSX4_A_F_Z_R,`ND3HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // ND3HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:29 and Version :1.1 //
 
//  START 
// CELL F_ND3HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_ND3HSX4_C_F_Z_R 0.1
`define F_ND3HSX4_C_R_Z_F 0.1
`define F_ND3HSX4_B_F_Z_R 0.1
`define F_ND3HSX4_B_R_Z_F 0.1
`define F_ND3HSX4_A_F_Z_R 0.1
`define F_ND3HSX4_A_R_Z_F 0.1

module F_ND3HSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C -=> Z) = (`F_ND3HSX4_C_F_Z_R,`F_ND3HSX4_C_R_Z_F);
      (B -=> Z) = (`F_ND3HSX4_B_F_Z_R,`F_ND3HSX4_B_R_Z_F);
      (A -=> Z) = (`F_ND3HSX4_A_F_Z_R,`F_ND3HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // F_ND3HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:29 and Version :1.1 //
 
//  START 
// CELL F_ND3HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_ND3HSX8_C_F_Z_R 0.1
`define F_ND3HSX8_C_R_Z_F 0.1
`define F_ND3HSX8_B_F_Z_R 0.1
`define F_ND3HSX8_B_R_Z_F 0.1
`define F_ND3HSX8_A_F_Z_R 0.1
`define F_ND3HSX8_A_R_Z_F 0.1

module F_ND3HSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C -=> Z) = (`F_ND3HSX8_C_F_Z_R,`F_ND3HSX8_C_R_Z_F);
      (B -=> Z) = (`F_ND3HSX8_B_F_Z_R,`F_ND3HSX8_B_R_Z_F);
      (A -=> Z) = (`F_ND3HSX8_A_F_Z_R,`F_ND3HSX8_A_R_Z_F);

   endspecify
`endif


endmodule // F_ND3HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:29 and Version :1.1 //
 
//  START 
// CELL M_ND3HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define M_ND3HSP_C_F_Z_R 0.1
`define M_ND3HSP_C_R_Z_F 0.1
`define M_ND3HSP_B_F_Z_R 0.1
`define M_ND3HSP_B_R_Z_F 0.1
`define M_ND3HSP_A_F_Z_R 0.1
`define M_ND3HSP_A_R_Z_F 0.1

module M_ND3HSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C -=> Z) = (`M_ND3HSP_C_F_Z_R,`M_ND3HSP_C_R_Z_F);
      (B -=> Z) = (`M_ND3HSP_B_F_Z_R,`M_ND3HSP_B_R_Z_F);
      (A -=> Z) = (`M_ND3HSP_A_F_Z_R,`M_ND3HSP_A_R_Z_F);

   endspecify
`endif


endmodule // M_ND3HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:29 and Version :1.1 //
 
//  START 
// CELL M_ND3HSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define M_ND3HSX3_C_F_Z_R 0.1
`define M_ND3HSX3_C_R_Z_F 0.1
`define M_ND3HSX3_B_F_Z_R 0.1
`define M_ND3HSX3_B_R_Z_F 0.1
`define M_ND3HSX3_A_F_Z_R 0.1
`define M_ND3HSX3_A_R_Z_F 0.1

module M_ND3HSX3 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C -=> Z) = (`M_ND3HSX3_C_F_Z_R,`M_ND3HSX3_C_R_Z_F);
      (B -=> Z) = (`M_ND3HSX3_B_F_Z_R,`M_ND3HSX3_B_R_Z_F);
      (A -=> Z) = (`M_ND3HSX3_A_F_Z_R,`M_ND3HSX3_A_R_Z_F);

   endspecify
`endif


endmodule // M_ND3HSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:29 and Version :1.1 //
 
//  START 
// CELL ND3AHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND3AHS_C_F_Z_R 0.1
`define ND3AHS_C_R_Z_F 0.1
`define ND3AHS_B_F_Z_R 0.1
`define ND3AHS_B_R_Z_F 0.1
`define ND3AHS_A_F_Z_F 0.1
`define ND3AHS_A_R_Z_R 0.1

module ND3AHS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`ND3AHS_C_F_Z_R,`ND3AHS_C_R_Z_F);
      (B -=> Z) = (`ND3AHS_B_F_Z_R,`ND3AHS_B_R_Z_F);
      (A +=> Z) = (`ND3AHS_A_R_Z_R,`ND3AHS_A_F_Z_F);

   endspecify
`endif


endmodule // ND3AHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:29 and Version :1.1 //
 
//  START 
// CELL ND3AHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND3AHSP_C_F_Z_R 0.1
`define ND3AHSP_C_R_Z_F 0.1
`define ND3AHSP_B_F_Z_R 0.1
`define ND3AHSP_B_R_Z_F 0.1
`define ND3AHSP_A_F_Z_F 0.1
`define ND3AHSP_A_R_Z_R 0.1

module ND3AHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`ND3AHSP_C_F_Z_R,`ND3AHSP_C_R_Z_F);
      (B -=> Z) = (`ND3AHSP_B_F_Z_R,`ND3AHSP_B_R_Z_F);
      (A +=> Z) = (`ND3AHSP_A_R_Z_R,`ND3AHSP_A_F_Z_F);

   endspecify
`endif


endmodule // ND3AHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:29 and Version :1.1 //
 
//  START 
// CELL ND3AHSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND3AHSX3_C_F_Z_R 0.1
`define ND3AHSX3_C_R_Z_F 0.1
`define ND3AHSX3_B_F_Z_R 0.1
`define ND3AHSX3_B_R_Z_F 0.1
`define ND3AHSX3_A_F_Z_F 0.1
`define ND3AHSX3_A_R_Z_R 0.1

module ND3AHSX3 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`ND3AHSX3_C_F_Z_R,`ND3AHSX3_C_R_Z_F);
      (B -=> Z) = (`ND3AHSX3_B_F_Z_R,`ND3AHSX3_B_R_Z_F);
      (A +=> Z) = (`ND3AHSX3_A_R_Z_R,`ND3AHSX3_A_F_Z_F);

   endspecify
`endif


endmodule // ND3AHSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:29 and Version :1.1 //
 
//  START 
// CELL ND3AHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND3AHSX4_C_F_Z_R 0.1
`define ND3AHSX4_C_R_Z_F 0.1
`define ND3AHSX4_B_F_Z_R 0.1
`define ND3AHSX4_B_R_Z_F 0.1
`define ND3AHSX4_A_F_Z_F 0.1
`define ND3AHSX4_A_R_Z_R 0.1

module ND3AHSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`ND3AHSX4_C_F_Z_R,`ND3AHSX4_C_R_Z_F);
      (B -=> Z) = (`ND3AHSX4_B_F_Z_R,`ND3AHSX4_B_R_Z_F);
      (A +=> Z) = (`ND3AHSX4_A_R_Z_R,`ND3AHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // ND3AHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:29 and Version :1.1 //
 
//  START 
// CELL F_ND3AHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_ND3AHSP_C_F_Z_R 0.1
`define F_ND3AHSP_C_R_Z_F 0.1
`define F_ND3AHSP_B_F_Z_R 0.1
`define F_ND3AHSP_B_R_Z_F 0.1
`define F_ND3AHSP_A_F_Z_F 0.1
`define F_ND3AHSP_A_R_Z_R 0.1

module F_ND3AHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`F_ND3AHSP_C_F_Z_R,`F_ND3AHSP_C_R_Z_F);
      (B -=> Z) = (`F_ND3AHSP_B_F_Z_R,`F_ND3AHSP_B_R_Z_F);
      (A +=> Z) = (`F_ND3AHSP_A_R_Z_R,`F_ND3AHSP_A_F_Z_F);

   endspecify
`endif


endmodule // F_ND3AHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:29 and Version :1.1 //
 
//  START 
// CELL F_ND3AHSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_ND3AHSX3_C_F_Z_R 0.1
`define F_ND3AHSX3_C_R_Z_F 0.1
`define F_ND3AHSX3_B_F_Z_R 0.1
`define F_ND3AHSX3_B_R_Z_F 0.1
`define F_ND3AHSX3_A_F_Z_F 0.1
`define F_ND3AHSX3_A_R_Z_R 0.1

module F_ND3AHSX3 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`F_ND3AHSX3_C_F_Z_R,`F_ND3AHSX3_C_R_Z_F);
      (B -=> Z) = (`F_ND3AHSX3_B_F_Z_R,`F_ND3AHSX3_B_R_Z_F);
      (A +=> Z) = (`F_ND3AHSX3_A_R_Z_R,`F_ND3AHSX3_A_F_Z_F);

   endspecify
`endif


endmodule // F_ND3AHSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:29 and Version :1.1 //
 
//  START 
// CELL F_ND3AHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_ND3AHSX4_C_F_Z_R 0.1
`define F_ND3AHSX4_C_R_Z_F 0.1
`define F_ND3AHSX4_B_F_Z_R 0.1
`define F_ND3AHSX4_B_R_Z_F 0.1
`define F_ND3AHSX4_A_F_Z_F 0.1
`define F_ND3AHSX4_A_R_Z_R 0.1

module F_ND3AHSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`F_ND3AHSX4_C_F_Z_R,`F_ND3AHSX4_C_R_Z_F);
      (B -=> Z) = (`F_ND3AHSX4_B_F_Z_R,`F_ND3AHSX4_B_R_Z_F);
      (A +=> Z) = (`F_ND3AHSX4_A_R_Z_R,`F_ND3AHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // F_ND3AHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:29 and Version :1.1 //
 
//  START 
// CELL F_ND3AHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_ND3AHSX8_C_F_Z_R 0.1
`define F_ND3AHSX8_C_R_Z_F 0.1
`define F_ND3AHSX8_B_F_Z_R 0.1
`define F_ND3AHSX8_B_R_Z_F 0.1
`define F_ND3AHSX8_A_F_Z_F 0.1
`define F_ND3AHSX8_A_R_Z_R 0.1

module F_ND3AHSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nand  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`F_ND3AHSX8_C_F_Z_R,`F_ND3AHSX8_C_R_Z_F);
      (B -=> Z) = (`F_ND3AHSX8_B_F_Z_R,`F_ND3AHSX8_B_R_Z_F);
      (A +=> Z) = (`F_ND3AHSX8_A_R_Z_R,`F_ND3AHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // F_ND3AHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:29 and Version :1.1 //
 
//  START 
// CELL ND4HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND4HSX05_D_F_Z_R 0.1
`define ND4HSX05_D_R_Z_F 0.1
`define ND4HSX05_C_F_Z_R 0.1
`define ND4HSX05_C_R_Z_F 0.1
`define ND4HSX05_B_F_Z_R 0.1
`define ND4HSX05_B_R_Z_F 0.1
`define ND4HSX05_A_F_Z_R 0.1
`define ND4HSX05_A_R_Z_F 0.1

module ND4HSX05 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`ND4HSX05_D_F_Z_R,`ND4HSX05_D_R_Z_F);
      (C -=> Z) = (`ND4HSX05_C_F_Z_R,`ND4HSX05_C_R_Z_F);
      (B -=> Z) = (`ND4HSX05_B_F_Z_R,`ND4HSX05_B_R_Z_F);
      (A -=> Z) = (`ND4HSX05_A_F_Z_R,`ND4HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // ND4HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:33 and Version :1.1 //
 
//  START 
// CELL ND4HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND4HS_D_F_Z_R 0.1
`define ND4HS_D_R_Z_F 0.1
`define ND4HS_C_F_Z_R 0.1
`define ND4HS_C_R_Z_F 0.1
`define ND4HS_B_F_Z_R 0.1
`define ND4HS_B_R_Z_F 0.1
`define ND4HS_A_F_Z_R 0.1
`define ND4HS_A_R_Z_F 0.1

module ND4HS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`ND4HS_D_F_Z_R,`ND4HS_D_R_Z_F);
      (C -=> Z) = (`ND4HS_C_F_Z_R,`ND4HS_C_R_Z_F);
      (B -=> Z) = (`ND4HS_B_F_Z_R,`ND4HS_B_R_Z_F);
      (A -=> Z) = (`ND4HS_A_F_Z_R,`ND4HS_A_R_Z_F);

   endspecify
`endif


endmodule // ND4HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:33 and Version :1.1 //
 
//  START 
// CELL ND4HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND4HSP_D_F_Z_R 0.1
`define ND4HSP_D_R_Z_F 0.1
`define ND4HSP_C_F_Z_R 0.1
`define ND4HSP_C_R_Z_F 0.1
`define ND4HSP_B_F_Z_R 0.1
`define ND4HSP_B_R_Z_F 0.1
`define ND4HSP_A_F_Z_R 0.1
`define ND4HSP_A_R_Z_F 0.1

module ND4HSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`ND4HSP_D_F_Z_R,`ND4HSP_D_R_Z_F);
      (C -=> Z) = (`ND4HSP_C_F_Z_R,`ND4HSP_C_R_Z_F);
      (B -=> Z) = (`ND4HSP_B_F_Z_R,`ND4HSP_B_R_Z_F);
      (A -=> Z) = (`ND4HSP_A_F_Z_R,`ND4HSP_A_R_Z_F);

   endspecify
`endif


endmodule // ND4HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:33 and Version :1.1 //
 
//  START 
// CELL ND4HSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND4HSX3_D_F_Z_R 0.1
`define ND4HSX3_D_R_Z_F 0.1
`define ND4HSX3_C_F_Z_R 0.1
`define ND4HSX3_C_R_Z_F 0.1
`define ND4HSX3_B_F_Z_R 0.1
`define ND4HSX3_B_R_Z_F 0.1
`define ND4HSX3_A_F_Z_R 0.1
`define ND4HSX3_A_R_Z_F 0.1

module ND4HSX3 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`ND4HSX3_D_F_Z_R,`ND4HSX3_D_R_Z_F);
      (C -=> Z) = (`ND4HSX3_C_F_Z_R,`ND4HSX3_C_R_Z_F);
      (B -=> Z) = (`ND4HSX3_B_F_Z_R,`ND4HSX3_B_R_Z_F);
      (A -=> Z) = (`ND4HSX3_A_F_Z_R,`ND4HSX3_A_R_Z_F);

   endspecify
`endif


endmodule // ND4HSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:33 and Version :1.1 //
 
//  START 
// CELL ND4HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND4HSX4_D_F_Z_R 0.1
`define ND4HSX4_D_R_Z_F 0.1
`define ND4HSX4_C_F_Z_R 0.1
`define ND4HSX4_C_R_Z_F 0.1
`define ND4HSX4_B_F_Z_R 0.1
`define ND4HSX4_B_R_Z_F 0.1
`define ND4HSX4_A_F_Z_R 0.1
`define ND4HSX4_A_R_Z_F 0.1

module ND4HSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`ND4HSX4_D_F_Z_R,`ND4HSX4_D_R_Z_F);
      (C -=> Z) = (`ND4HSX4_C_F_Z_R,`ND4HSX4_C_R_Z_F);
      (B -=> Z) = (`ND4HSX4_B_F_Z_R,`ND4HSX4_B_R_Z_F);
      (A -=> Z) = (`ND4HSX4_A_F_Z_R,`ND4HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // ND4HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:33 and Version :1.1 //
 
//  START 
// CELL F_ND4HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_ND4HS_D_F_Z_R 0.1
`define F_ND4HS_D_R_Z_F 0.1
`define F_ND4HS_C_F_Z_R 0.1
`define F_ND4HS_C_R_Z_F 0.1
`define F_ND4HS_B_F_Z_R 0.1
`define F_ND4HS_B_R_Z_F 0.1
`define F_ND4HS_A_F_Z_R 0.1
`define F_ND4HS_A_R_Z_F 0.1

module F_ND4HS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`F_ND4HS_D_F_Z_R,`F_ND4HS_D_R_Z_F);
      (C -=> Z) = (`F_ND4HS_C_F_Z_R,`F_ND4HS_C_R_Z_F);
      (B -=> Z) = (`F_ND4HS_B_F_Z_R,`F_ND4HS_B_R_Z_F);
      (A -=> Z) = (`F_ND4HS_A_F_Z_R,`F_ND4HS_A_R_Z_F);

   endspecify
`endif


endmodule // F_ND4HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:33 and Version :1.1 //
 
//  START 
// CELL F_ND4HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_ND4HSP_D_F_Z_R 0.1
`define F_ND4HSP_D_R_Z_F 0.1
`define F_ND4HSP_C_F_Z_R 0.1
`define F_ND4HSP_C_R_Z_F 0.1
`define F_ND4HSP_B_F_Z_R 0.1
`define F_ND4HSP_B_R_Z_F 0.1
`define F_ND4HSP_A_F_Z_R 0.1
`define F_ND4HSP_A_R_Z_F 0.1

module F_ND4HSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`F_ND4HSP_D_F_Z_R,`F_ND4HSP_D_R_Z_F);
      (C -=> Z) = (`F_ND4HSP_C_F_Z_R,`F_ND4HSP_C_R_Z_F);
      (B -=> Z) = (`F_ND4HSP_B_F_Z_R,`F_ND4HSP_B_R_Z_F);
      (A -=> Z) = (`F_ND4HSP_A_F_Z_R,`F_ND4HSP_A_R_Z_F);

   endspecify
`endif


endmodule // F_ND4HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:33 and Version :1.1 //
 
//  START 
// CELL ND4HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND4HSX8_D_F_Z_R 0.1
`define ND4HSX8_D_R_Z_F 0.1
`define ND4HSX8_C_F_Z_R 0.1
`define ND4HSX8_C_R_Z_F 0.1
`define ND4HSX8_B_F_Z_R 0.1
`define ND4HSX8_B_R_Z_F 0.1
`define ND4HSX8_A_F_Z_R 0.1
`define ND4HSX8_A_R_Z_F 0.1

module ND4HSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nand  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`ND4HSX8_D_F_Z_R,`ND4HSX8_D_R_Z_F);
      (C -=> Z) = (`ND4HSX8_C_F_Z_R,`ND4HSX8_C_R_Z_F);
      (B -=> Z) = (`ND4HSX8_B_F_Z_R,`ND4HSX8_B_R_Z_F);
      (A -=> Z) = (`ND4HSX8_A_F_Z_R,`ND4HSX8_A_R_Z_F);

   endspecify
`endif


endmodule // ND4HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:33 and Version :1.1 //
 
//  START 
// CELL ND5HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND5HS_E_F_Z_R 0.1
`define ND5HS_E_R_Z_F 0.1
`define ND5HS_D_F_Z_R 0.1
`define ND5HS_D_R_Z_F 0.1
`define ND5HS_C_F_Z_R 0.1
`define ND5HS_C_R_Z_F 0.1
`define ND5HS_B_F_Z_R 0.1
`define ND5HS_B_R_Z_F 0.1
`define ND5HS_A_F_Z_R 0.1
`define ND5HS_A_R_Z_F 0.1

module ND5HS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   nand  u0 (Z, A, B, C, D, E);


`ifdef functional
`else
   specify

      (E -=> Z) = (`ND5HS_E_F_Z_R,`ND5HS_E_R_Z_F);
      (D -=> Z) = (`ND5HS_D_F_Z_R,`ND5HS_D_R_Z_F);
      (C -=> Z) = (`ND5HS_C_F_Z_R,`ND5HS_C_R_Z_F);
      (B -=> Z) = (`ND5HS_B_F_Z_R,`ND5HS_B_R_Z_F);
      (A -=> Z) = (`ND5HS_A_F_Z_R,`ND5HS_A_R_Z_F);

   endspecify
`endif


endmodule // ND5HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:40 and Version :1.1 //
 
//  START 
// CELL ND5HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND5HSP_E_F_Z_R 0.1
`define ND5HSP_E_R_Z_F 0.1
`define ND5HSP_D_F_Z_R 0.1
`define ND5HSP_D_R_Z_F 0.1
`define ND5HSP_C_F_Z_R 0.1
`define ND5HSP_C_R_Z_F 0.1
`define ND5HSP_B_F_Z_R 0.1
`define ND5HSP_B_R_Z_F 0.1
`define ND5HSP_A_F_Z_R 0.1
`define ND5HSP_A_R_Z_F 0.1

module ND5HSP (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   nand  u0 (Z, A, B, C, D, E);


`ifdef functional
`else
   specify

      (E -=> Z) = (`ND5HSP_E_F_Z_R,`ND5HSP_E_R_Z_F);
      (D -=> Z) = (`ND5HSP_D_F_Z_R,`ND5HSP_D_R_Z_F);
      (C -=> Z) = (`ND5HSP_C_F_Z_R,`ND5HSP_C_R_Z_F);
      (B -=> Z) = (`ND5HSP_B_F_Z_R,`ND5HSP_B_R_Z_F);
      (A -=> Z) = (`ND5HSP_A_F_Z_R,`ND5HSP_A_R_Z_F);

   endspecify
`endif


endmodule // ND5HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:40 and Version :1.1 //
 
//  START 
// CELL ND5HSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND5HSX3_E_F_Z_R 0.1
`define ND5HSX3_E_R_Z_F 0.1
`define ND5HSX3_D_F_Z_R 0.1
`define ND5HSX3_D_R_Z_F 0.1
`define ND5HSX3_C_F_Z_R 0.1
`define ND5HSX3_C_R_Z_F 0.1
`define ND5HSX3_B_F_Z_R 0.1
`define ND5HSX3_B_R_Z_F 0.1
`define ND5HSX3_A_F_Z_R 0.1
`define ND5HSX3_A_R_Z_F 0.1

module ND5HSX3 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   nand  u0 (Z, A, B, C, D, E);


`ifdef functional
`else
   specify

      (E -=> Z) = (`ND5HSX3_E_F_Z_R,`ND5HSX3_E_R_Z_F);
      (D -=> Z) = (`ND5HSX3_D_F_Z_R,`ND5HSX3_D_R_Z_F);
      (C -=> Z) = (`ND5HSX3_C_F_Z_R,`ND5HSX3_C_R_Z_F);
      (B -=> Z) = (`ND5HSX3_B_F_Z_R,`ND5HSX3_B_R_Z_F);
      (A -=> Z) = (`ND5HSX3_A_F_Z_R,`ND5HSX3_A_R_Z_F);

   endspecify
`endif


endmodule // ND5HSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:40 and Version :1.1 //
 
//  START 
// CELL ND5HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND5HSX4_E_F_Z_R 0.1
`define ND5HSX4_E_R_Z_F 0.1
`define ND5HSX4_D_F_Z_R 0.1
`define ND5HSX4_D_R_Z_F 0.1
`define ND5HSX4_C_F_Z_R 0.1
`define ND5HSX4_C_R_Z_F 0.1
`define ND5HSX4_B_F_Z_R 0.1
`define ND5HSX4_B_R_Z_F 0.1
`define ND5HSX4_A_F_Z_R 0.1
`define ND5HSX4_A_R_Z_F 0.1

module ND5HSX4 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   nand  u0 (Z, A, B, C, D, E);


`ifdef functional
`else
   specify

      (E -=> Z) = (`ND5HSX4_E_F_Z_R,`ND5HSX4_E_R_Z_F);
      (D -=> Z) = (`ND5HSX4_D_F_Z_R,`ND5HSX4_D_R_Z_F);
      (C -=> Z) = (`ND5HSX4_C_F_Z_R,`ND5HSX4_C_R_Z_F);
      (B -=> Z) = (`ND5HSX4_B_F_Z_R,`ND5HSX4_B_R_Z_F);
      (A -=> Z) = (`ND5HSX4_A_F_Z_R,`ND5HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // ND5HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:40 and Version :1.1 //
 
//  START 
// CELL ND6HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND6HS_F_F_Z_R 0.1
`define ND6HS_F_R_Z_F 0.1
`define ND6HS_E_F_Z_R 0.1
`define ND6HS_E_R_Z_F 0.1
`define ND6HS_D_F_Z_R 0.1
`define ND6HS_D_R_Z_F 0.1
`define ND6HS_C_F_Z_R 0.1
`define ND6HS_C_R_Z_F 0.1
`define ND6HS_B_F_Z_R 0.1
`define ND6HS_B_R_Z_F 0.1
`define ND6HS_A_F_Z_R 0.1
`define ND6HS_A_R_Z_F 0.1

module ND6HS (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   nand  u0 (Z, A, B, C, D, E, F);


`ifdef functional
`else
   specify

      (F -=> Z) = (`ND6HS_F_F_Z_R,`ND6HS_F_R_Z_F);
      (E -=> Z) = (`ND6HS_E_F_Z_R,`ND6HS_E_R_Z_F);
      (D -=> Z) = (`ND6HS_D_F_Z_R,`ND6HS_D_R_Z_F);
      (C -=> Z) = (`ND6HS_C_F_Z_R,`ND6HS_C_R_Z_F);
      (B -=> Z) = (`ND6HS_B_F_Z_R,`ND6HS_B_R_Z_F);
      (A -=> Z) = (`ND6HS_A_F_Z_R,`ND6HS_A_R_Z_F);

   endspecify
`endif


endmodule // ND6HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:43 and Version :1.1 //
 
//  START 
// CELL ND6HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND6HSP_F_F_Z_R 0.1
`define ND6HSP_F_R_Z_F 0.1
`define ND6HSP_E_F_Z_R 0.1
`define ND6HSP_E_R_Z_F 0.1
`define ND6HSP_D_F_Z_R 0.1
`define ND6HSP_D_R_Z_F 0.1
`define ND6HSP_C_F_Z_R 0.1
`define ND6HSP_C_R_Z_F 0.1
`define ND6HSP_B_F_Z_R 0.1
`define ND6HSP_B_R_Z_F 0.1
`define ND6HSP_A_F_Z_R 0.1
`define ND6HSP_A_R_Z_F 0.1

module ND6HSP (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   nand  u0 (Z, A, B, C, D, E, F);


`ifdef functional
`else
   specify

      (F -=> Z) = (`ND6HSP_F_F_Z_R,`ND6HSP_F_R_Z_F);
      (E -=> Z) = (`ND6HSP_E_F_Z_R,`ND6HSP_E_R_Z_F);
      (D -=> Z) = (`ND6HSP_D_F_Z_R,`ND6HSP_D_R_Z_F);
      (C -=> Z) = (`ND6HSP_C_F_Z_R,`ND6HSP_C_R_Z_F);
      (B -=> Z) = (`ND6HSP_B_F_Z_R,`ND6HSP_B_R_Z_F);
      (A -=> Z) = (`ND6HSP_A_F_Z_R,`ND6HSP_A_R_Z_F);

   endspecify
`endif


endmodule // ND6HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:43 and Version :1.1 //
 
//  START 
// CELL ND7HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND7HS_G_F_Z_R 0.1
`define ND7HS_G_R_Z_F 0.1
`define ND7HS_F_F_Z_R 0.1
`define ND7HS_F_R_Z_F 0.1
`define ND7HS_E_F_Z_R 0.1
`define ND7HS_E_R_Z_F 0.1
`define ND7HS_D_F_Z_R 0.1
`define ND7HS_D_R_Z_F 0.1
`define ND7HS_C_F_Z_R 0.1
`define ND7HS_C_R_Z_F 0.1
`define ND7HS_B_F_Z_R 0.1
`define ND7HS_B_R_Z_F 0.1
`define ND7HS_A_F_Z_R 0.1
`define ND7HS_A_R_Z_F 0.1

module ND7HS (Z, A, B, C, D, E, F, G);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;
   input G;


   nand  u0 (Z, A, B, C, D, E, F, G);


`ifdef functional
`else
   specify

      (G -=> Z) = (`ND7HS_G_F_Z_R,`ND7HS_G_R_Z_F);
      (F -=> Z) = (`ND7HS_F_F_Z_R,`ND7HS_F_R_Z_F);
      (E -=> Z) = (`ND7HS_E_F_Z_R,`ND7HS_E_R_Z_F);
      (D -=> Z) = (`ND7HS_D_F_Z_R,`ND7HS_D_R_Z_F);
      (C -=> Z) = (`ND7HS_C_F_Z_R,`ND7HS_C_R_Z_F);
      (B -=> Z) = (`ND7HS_B_F_Z_R,`ND7HS_B_R_Z_F);
      (A -=> Z) = (`ND7HS_A_F_Z_R,`ND7HS_A_R_Z_F);

   endspecify
`endif


endmodule // ND7HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:50 and Version :1.1 //
 
//  START 
// CELL ND8HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND8HS_H_F_Z_R 0.1
`define ND8HS_H_R_Z_F 0.1
`define ND8HS_G_F_Z_R 0.1
`define ND8HS_G_R_Z_F 0.1
`define ND8HS_F_F_Z_R 0.1
`define ND8HS_F_R_Z_F 0.1
`define ND8HS_E_F_Z_R 0.1
`define ND8HS_E_R_Z_F 0.1
`define ND8HS_D_F_Z_R 0.1
`define ND8HS_D_R_Z_F 0.1
`define ND8HS_C_F_Z_R 0.1
`define ND8HS_C_R_Z_F 0.1
`define ND8HS_B_F_Z_R 0.1
`define ND8HS_B_R_Z_F 0.1
`define ND8HS_A_F_Z_R 0.1
`define ND8HS_A_R_Z_F 0.1

module ND8HS (Z, A, B, C, D, E, F, G, H);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;
   input G;
   input H;


   nand  u0 (Z, A, B, C, D, E, F, G, H);


`ifdef functional
`else
   specify

      (H -=> Z) = (`ND8HS_H_F_Z_R,`ND8HS_H_R_Z_F);
      (G -=> Z) = (`ND8HS_G_F_Z_R,`ND8HS_G_R_Z_F);
      (F -=> Z) = (`ND8HS_F_F_Z_R,`ND8HS_F_R_Z_F);
      (E -=> Z) = (`ND8HS_E_F_Z_R,`ND8HS_E_R_Z_F);
      (D -=> Z) = (`ND8HS_D_F_Z_R,`ND8HS_D_R_Z_F);
      (C -=> Z) = (`ND8HS_C_F_Z_R,`ND8HS_C_R_Z_F);
      (B -=> Z) = (`ND8HS_B_F_Z_R,`ND8HS_B_R_Z_F);
      (A -=> Z) = (`ND8HS_A_F_Z_R,`ND8HS_A_R_Z_F);

   endspecify
`endif


endmodule // ND8HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:50 and Version :1.1 //
 
//  START 
// CELL ND8HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define ND8HSP_H_F_Z_R 0.1
`define ND8HSP_H_R_Z_F 0.1
`define ND8HSP_G_F_Z_R 0.1
`define ND8HSP_G_R_Z_F 0.1
`define ND8HSP_F_F_Z_R 0.1
`define ND8HSP_F_R_Z_F 0.1
`define ND8HSP_E_F_Z_R 0.1
`define ND8HSP_E_R_Z_F 0.1
`define ND8HSP_D_F_Z_R 0.1
`define ND8HSP_D_R_Z_F 0.1
`define ND8HSP_C_F_Z_R 0.1
`define ND8HSP_C_R_Z_F 0.1
`define ND8HSP_B_F_Z_R 0.1
`define ND8HSP_B_R_Z_F 0.1
`define ND8HSP_A_F_Z_R 0.1
`define ND8HSP_A_R_Z_F 0.1

module ND8HSP (Z, A, B, C, D, E, F, G, H);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;
   input G;
   input H;


   nand  u0 (Z, A, B, C, D, E, F, G, H);


`ifdef functional
`else
   specify

      (H -=> Z) = (`ND8HSP_H_F_Z_R,`ND8HSP_H_R_Z_F);
      (G -=> Z) = (`ND8HSP_G_F_Z_R,`ND8HSP_G_R_Z_F);
      (F -=> Z) = (`ND8HSP_F_F_Z_R,`ND8HSP_F_R_Z_F);
      (E -=> Z) = (`ND8HSP_E_F_Z_R,`ND8HSP_E_R_Z_F);
      (D -=> Z) = (`ND8HSP_D_F_Z_R,`ND8HSP_D_R_Z_F);
      (C -=> Z) = (`ND8HSP_C_F_Z_R,`ND8HSP_C_R_Z_F);
      (B -=> Z) = (`ND8HSP_B_F_Z_R,`ND8HSP_B_R_Z_F);
      (A -=> Z) = (`ND8HSP_A_F_Z_R,`ND8HSP_A_R_Z_F);

   endspecify
`endif


endmodule // ND8HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:50 and Version :1.1 //
 
//  START 
// CELL NR2HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR2HSX05_B_F_Z_R 0.1
`define NR2HSX05_B_R_Z_F 0.1
`define NR2HSX05_A_F_Z_R 0.1
`define NR2HSX05_A_R_Z_F 0.1

module NR2HSX05 (Z, A, B);

   output Z;
   input A;
   input B;


   nor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`NR2HSX05_B_F_Z_R,`NR2HSX05_B_R_Z_F);
      (A -=> Z) = (`NR2HSX05_A_F_Z_R,`NR2HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // NR2HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START 
// CELL NR2HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR2HS_B_F_Z_R 0.1
`define NR2HS_B_R_Z_F 0.1
`define NR2HS_A_F_Z_R 0.1
`define NR2HS_A_R_Z_F 0.1

module NR2HS (Z, A, B);

   output Z;
   input A;
   input B;


   nor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`NR2HS_B_F_Z_R,`NR2HS_B_R_Z_F);
      (A -=> Z) = (`NR2HS_A_F_Z_R,`NR2HS_A_R_Z_F);

   endspecify
`endif


endmodule // NR2HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START 
// CELL NR2HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR2HSP_B_F_Z_R 0.1
`define NR2HSP_B_R_Z_F 0.1
`define NR2HSP_A_F_Z_R 0.1
`define NR2HSP_A_R_Z_F 0.1

module NR2HSP (Z, A, B);

   output Z;
   input A;
   input B;


   nor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`NR2HSP_B_F_Z_R,`NR2HSP_B_R_Z_F);
      (A -=> Z) = (`NR2HSP_A_F_Z_R,`NR2HSP_A_R_Z_F);

   endspecify
`endif


endmodule // NR2HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START 
// CELL NR2HSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR2HSX3_B_F_Z_R 0.1
`define NR2HSX3_B_R_Z_F 0.1
`define NR2HSX3_A_F_Z_R 0.1
`define NR2HSX3_A_R_Z_F 0.1

module NR2HSX3 (Z, A, B);

   output Z;
   input A;
   input B;


   nor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`NR2HSX3_B_F_Z_R,`NR2HSX3_B_R_Z_F);
      (A -=> Z) = (`NR2HSX3_A_F_Z_R,`NR2HSX3_A_R_Z_F);

   endspecify
`endif


endmodule // NR2HSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START 
// CELL NR2HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR2HSX4_B_F_Z_R 0.1
`define NR2HSX4_B_R_Z_F 0.1
`define NR2HSX4_A_F_Z_R 0.1
`define NR2HSX4_A_R_Z_F 0.1

module NR2HSX4 (Z, A, B);

   output Z;
   input A;
   input B;


   nor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`NR2HSX4_B_F_Z_R,`NR2HSX4_B_R_Z_F);
      (A -=> Z) = (`NR2HSX4_A_F_Z_R,`NR2HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // NR2HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START 
// CELL F_NR2HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_NR2HSP_B_F_Z_R 0.1
`define F_NR2HSP_B_R_Z_F 0.1
`define F_NR2HSP_A_F_Z_R 0.1
`define F_NR2HSP_A_R_Z_F 0.1

module F_NR2HSP (Z, A, B);

   output Z;
   input A;
   input B;


   nor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`F_NR2HSP_B_F_Z_R,`F_NR2HSP_B_R_Z_F);
      (A -=> Z) = (`F_NR2HSP_A_F_Z_R,`F_NR2HSP_A_R_Z_F);

   endspecify
`endif


endmodule // F_NR2HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START 
// CELL F_NR2HSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_NR2HSX3_B_F_Z_R 0.1
`define F_NR2HSX3_B_R_Z_F 0.1
`define F_NR2HSX3_A_F_Z_R 0.1
`define F_NR2HSX3_A_R_Z_F 0.1

module F_NR2HSX3 (Z, A, B);

   output Z;
   input A;
   input B;


   nor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`F_NR2HSX3_B_F_Z_R,`F_NR2HSX3_B_R_Z_F);
      (A -=> Z) = (`F_NR2HSX3_A_F_Z_R,`F_NR2HSX3_A_R_Z_F);

   endspecify
`endif


endmodule // F_NR2HSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START 
// CELL F_NR2HSX6

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_NR2HSX6_B_F_Z_R 0.1
`define F_NR2HSX6_B_R_Z_F 0.1
`define F_NR2HSX6_A_F_Z_R 0.1
`define F_NR2HSX6_A_R_Z_F 0.1

module F_NR2HSX6 (Z, A, B);

   output Z;
   input A;
   input B;


   nor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`F_NR2HSX6_B_F_Z_R,`F_NR2HSX6_B_R_Z_F);
      (A -=> Z) = (`F_NR2HSX6_A_F_Z_R,`F_NR2HSX6_A_R_Z_F);

   endspecify
`endif


endmodule // F_NR2HSX6
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START 
// CELL M_NR2HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define M_NR2HS_B_F_Z_R 0.1
`define M_NR2HS_B_R_Z_F 0.1
`define M_NR2HS_A_F_Z_R 0.1
`define M_NR2HS_A_R_Z_F 0.1

module M_NR2HS (Z, A, B);

   output Z;
   input A;
   input B;


   nor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`M_NR2HS_B_F_Z_R,`M_NR2HS_B_R_Z_F);
      (A -=> Z) = (`M_NR2HS_A_F_Z_R,`M_NR2HS_A_R_Z_F);

   endspecify
`endif


endmodule // M_NR2HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START 
// CELL NR2HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR2HSX8_B_F_Z_R 0.1
`define NR2HSX8_B_R_Z_F 0.1
`define NR2HSX8_A_F_Z_R 0.1
`define NR2HSX8_A_R_Z_F 0.1

module NR2HSX8 (Z, A, B);

   output Z;
   input A;
   input B;


   nor  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`NR2HSX8_B_F_Z_R,`NR2HSX8_B_R_Z_F);
      (A -=> Z) = (`NR2HSX8_A_F_Z_R,`NR2HSX8_A_R_Z_F);

   endspecify
`endif


endmodule // NR2HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START 
// CELL NR2AHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR2AHS_B_F_Z_R 0.1
`define NR2AHS_B_R_Z_F 0.1
`define NR2AHS_A_F_Z_F 0.1
`define NR2AHS_A_R_Z_R 0.1

module NR2AHS (Z, A, B);

   output Z;
   input A;
   input B;


   and  u0 (Z, A, BX);
   not  u1 (BX, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`NR2AHS_B_F_Z_R,`NR2AHS_B_R_Z_F);
      (A +=> Z) = (`NR2AHS_A_R_Z_R,`NR2AHS_A_F_Z_F);

   endspecify
`endif


endmodule // NR2AHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START 
// CELL NR2AHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR2AHSP_B_F_Z_R 0.1
`define NR2AHSP_B_R_Z_F 0.1
`define NR2AHSP_A_F_Z_F 0.1
`define NR2AHSP_A_R_Z_R 0.1

module NR2AHSP (Z, A, B);

   output Z;
   input A;
   input B;


   and  u0 (Z, A, BX);
   not  u1 (BX, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`NR2AHSP_B_F_Z_R,`NR2AHSP_B_R_Z_F);
      (A +=> Z) = (`NR2AHSP_A_R_Z_R,`NR2AHSP_A_F_Z_F);

   endspecify
`endif


endmodule // NR2AHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START 
// CELL NR2AHSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR2AHSX3_B_F_Z_R 0.1
`define NR2AHSX3_B_R_Z_F 0.1
`define NR2AHSX3_A_F_Z_F 0.1
`define NR2AHSX3_A_R_Z_R 0.1

module NR2AHSX3 (Z, A, B);

   output Z;
   input A;
   input B;


   and  u0 (Z, A, BX);
   not  u1 (BX, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`NR2AHSX3_B_F_Z_R,`NR2AHSX3_B_R_Z_F);
      (A +=> Z) = (`NR2AHSX3_A_R_Z_R,`NR2AHSX3_A_F_Z_F);

   endspecify
`endif


endmodule // NR2AHSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START 
// CELL NR2AHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR2AHSX4_B_F_Z_R 0.1
`define NR2AHSX4_B_R_Z_F 0.1
`define NR2AHSX4_A_F_Z_F 0.1
`define NR2AHSX4_A_R_Z_R 0.1

module NR2AHSX4 (Z, A, B);

   output Z;
   input A;
   input B;


   and  u0 (Z, A, BX);
   not  u1 (BX, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`NR2AHSX4_B_F_Z_R,`NR2AHSX4_B_R_Z_F);
      (A +=> Z) = (`NR2AHSX4_A_R_Z_R,`NR2AHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // NR2AHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START 
// CELL F_NR2AHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_NR2AHSP_B_F_Z_R 0.1
`define F_NR2AHSP_B_R_Z_F 0.1
`define F_NR2AHSP_A_F_Z_F 0.1
`define F_NR2AHSP_A_R_Z_R 0.1

module F_NR2AHSP (Z, A, B);

   output Z;
   input A;
   input B;


   and  u0 (Z, A, BX);
   not  u1 (BX, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`F_NR2AHSP_B_F_Z_R,`F_NR2AHSP_B_R_Z_F);
      (A +=> Z) = (`F_NR2AHSP_A_R_Z_R,`F_NR2AHSP_A_F_Z_F);

   endspecify
`endif


endmodule // F_NR2AHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START 
// CELL F_NR2AHSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_NR2AHSX3_B_F_Z_R 0.1
`define F_NR2AHSX3_B_R_Z_F 0.1
`define F_NR2AHSX3_A_F_Z_F 0.1
`define F_NR2AHSX3_A_R_Z_R 0.1

module F_NR2AHSX3 (Z, A, B);

   output Z;
   input A;
   input B;


   and  u0 (Z, A, BX);
   not  u1 (BX, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`F_NR2AHSX3_B_F_Z_R,`F_NR2AHSX3_B_R_Z_F);
      (A +=> Z) = (`F_NR2AHSX3_A_R_Z_R,`F_NR2AHSX3_A_F_Z_F);

   endspecify
`endif


endmodule // F_NR2AHSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START 
// CELL NR2AHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR2AHSX8_B_F_Z_R 0.1
`define NR2AHSX8_B_R_Z_F 0.1
`define NR2AHSX8_A_F_Z_F 0.1
`define NR2AHSX8_A_R_Z_R 0.1

module NR2AHSX8 (Z, A, B);

   output Z;
   input A;
   input B;


   and  u0 (Z, A, BX);
   not  u1 (BX, B);


`ifdef functional
`else
   specify

      (B -=> Z) = (`NR2AHSX8_B_F_Z_R,`NR2AHSX8_B_R_Z_F);
      (A +=> Z) = (`NR2AHSX8_A_R_Z_R,`NR2AHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // NR2AHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:57 and Version :1.1 //
 
//  START 
// CELL NR3HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR3HSX05_C_F_Z_R 0.1
`define NR3HSX05_C_R_Z_F 0.1
`define NR3HSX05_B_F_Z_R 0.1
`define NR3HSX05_B_R_Z_F 0.1
`define NR3HSX05_A_F_Z_R 0.1
`define NR3HSX05_A_R_Z_F 0.1

module NR3HSX05 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C -=> Z) = (`NR3HSX05_C_F_Z_R,`NR3HSX05_C_R_Z_F);
      (B -=> Z) = (`NR3HSX05_B_F_Z_R,`NR3HSX05_B_R_Z_F);
      (A -=> Z) = (`NR3HSX05_A_F_Z_R,`NR3HSX05_A_R_Z_F);

   endspecify
`endif


endmodule
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:59 and Version :1.1 //
 
//  START 
// CELL NR3HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR3HS_C_F_Z_R 0.1
`define NR3HS_C_R_Z_F 0.1
`define NR3HS_B_F_Z_R 0.1
`define NR3HS_B_R_Z_F 0.1
`define NR3HS_A_F_Z_R 0.1
`define NR3HS_A_R_Z_F 0.1

module NR3HS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C -=> Z) = (`NR3HS_C_F_Z_R,`NR3HS_C_R_Z_F);
      (B -=> Z) = (`NR3HS_B_F_Z_R,`NR3HS_B_R_Z_F);
      (A -=> Z) = (`NR3HS_A_F_Z_R,`NR3HS_A_R_Z_F);

   endspecify
`endif


endmodule
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:59 and Version :1.1 //
 
//  START 
// CELL NR3HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR3HSP_C_F_Z_R 0.1
`define NR3HSP_C_R_Z_F 0.1
`define NR3HSP_B_F_Z_R 0.1
`define NR3HSP_B_R_Z_F 0.1
`define NR3HSP_A_F_Z_R 0.1
`define NR3HSP_A_R_Z_F 0.1

module NR3HSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C -=> Z) = (`NR3HSP_C_F_Z_R,`NR3HSP_C_R_Z_F);
      (B -=> Z) = (`NR3HSP_B_F_Z_R,`NR3HSP_B_R_Z_F);
      (A -=> Z) = (`NR3HSP_A_F_Z_R,`NR3HSP_A_R_Z_F);

   endspecify
`endif


endmodule
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:59 and Version :1.1 //
 
//  START 
// CELL NR3HSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR3HSX3_C_F_Z_R 0.1
`define NR3HSX3_C_R_Z_F 0.1
`define NR3HSX3_B_F_Z_R 0.1
`define NR3HSX3_B_R_Z_F 0.1
`define NR3HSX3_A_F_Z_R 0.1
`define NR3HSX3_A_R_Z_F 0.1

module NR3HSX3 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C -=> Z) = (`NR3HSX3_C_F_Z_R,`NR3HSX3_C_R_Z_F);
      (B -=> Z) = (`NR3HSX3_B_F_Z_R,`NR3HSX3_B_R_Z_F);
      (A -=> Z) = (`NR3HSX3_A_F_Z_R,`NR3HSX3_A_R_Z_F);

   endspecify
`endif


endmodule
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:59 and Version :1.1 //
 
//  START 
// CELL NR3HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR3HSX4_C_F_Z_R 0.1
`define NR3HSX4_C_R_Z_F 0.1
`define NR3HSX4_B_F_Z_R 0.1
`define NR3HSX4_B_R_Z_F 0.1
`define NR3HSX4_A_F_Z_R 0.1
`define NR3HSX4_A_R_Z_F 0.1

module NR3HSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C -=> Z) = (`NR3HSX4_C_F_Z_R,`NR3HSX4_C_R_Z_F);
      (B -=> Z) = (`NR3HSX4_B_F_Z_R,`NR3HSX4_B_R_Z_F);
      (A -=> Z) = (`NR3HSX4_A_F_Z_R,`NR3HSX4_A_R_Z_F);

   endspecify
`endif


endmodule
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:59 and Version :1.1 //
 
//  START 
// CELL F_NR3HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_NR3HS_C_F_Z_R 0.1
`define F_NR3HS_C_R_Z_F 0.1
`define F_NR3HS_B_F_Z_R 0.1
`define F_NR3HS_B_R_Z_F 0.1
`define F_NR3HS_A_F_Z_R 0.1
`define F_NR3HS_A_R_Z_F 0.1

module F_NR3HS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C -=> Z) = (`F_NR3HS_C_F_Z_R,`F_NR3HS_C_R_Z_F);
      (B -=> Z) = (`F_NR3HS_B_F_Z_R,`F_NR3HS_B_R_Z_F);
      (A -=> Z) = (`F_NR3HS_A_F_Z_R,`F_NR3HS_A_R_Z_F);

   endspecify
`endif


endmodule
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:59 and Version :1.1 //
 
//  START 
// CELL F_NR3HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_NR3HSP_C_F_Z_R 0.1
`define F_NR3HSP_C_R_Z_F 0.1
`define F_NR3HSP_B_F_Z_R 0.1
`define F_NR3HSP_B_R_Z_F 0.1
`define F_NR3HSP_A_F_Z_R 0.1
`define F_NR3HSP_A_R_Z_F 0.1

module F_NR3HSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C -=> Z) = (`F_NR3HSP_C_F_Z_R,`F_NR3HSP_C_R_Z_F);
      (B -=> Z) = (`F_NR3HSP_B_F_Z_R,`F_NR3HSP_B_R_Z_F);
      (A -=> Z) = (`F_NR3HSP_A_F_Z_R,`F_NR3HSP_A_R_Z_F);

   endspecify
`endif


endmodule
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:59 and Version :1.1 //
 
//  START 
// CELL NR3HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR3HSX8_C_F_Z_R 0.1
`define NR3HSX8_C_R_Z_F 0.1
`define NR3HSX8_B_F_Z_R 0.1
`define NR3HSX8_B_R_Z_F 0.1
`define NR3HSX8_A_F_Z_R 0.1
`define NR3HSX8_A_R_Z_F 0.1

module NR3HSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C -=> Z) = (`NR3HSX8_C_F_Z_R,`NR3HSX8_C_R_Z_F);
      (B -=> Z) = (`NR3HSX8_B_F_Z_R,`NR3HSX8_B_R_Z_F);
      (A -=> Z) = (`NR3HSX8_A_F_Z_R,`NR3HSX8_A_R_Z_F);

   endspecify
`endif


endmodule
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:19:59 and Version :1.1 //
 
//  START 
// CELL NR3AHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR3AHS_C_F_Z_R 0.1
`define NR3AHS_C_R_Z_F 0.1
`define NR3AHS_B_F_Z_R 0.1
`define NR3AHS_B_R_Z_F 0.1
`define NR3AHS_A_F_Z_F 0.1
`define NR3AHS_A_R_Z_R 0.1

module NR3AHS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`NR3AHS_C_F_Z_R,`NR3AHS_C_R_Z_F);
      (B -=> Z) = (`NR3AHS_B_F_Z_R,`NR3AHS_B_R_Z_F);
      (A +=> Z) = (`NR3AHS_A_R_Z_R,`NR3AHS_A_F_Z_F);

   endspecify
`endif


endmodule // NR3AHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:03 and Version :1.1 //
 
//  START 
// CELL NR3AHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR3AHSP_C_F_Z_R 0.1
`define NR3AHSP_C_R_Z_F 0.1
`define NR3AHSP_B_F_Z_R 0.1
`define NR3AHSP_B_R_Z_F 0.1
`define NR3AHSP_A_F_Z_F 0.1
`define NR3AHSP_A_R_Z_R 0.1

module NR3AHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`NR3AHSP_C_F_Z_R,`NR3AHSP_C_R_Z_F);
      (B -=> Z) = (`NR3AHSP_B_F_Z_R,`NR3AHSP_B_R_Z_F);
      (A +=> Z) = (`NR3AHSP_A_R_Z_R,`NR3AHSP_A_F_Z_F);

   endspecify
`endif


endmodule // NR3AHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:03 and Version :1.1 //
 
//  START 
// CELL NR3AHSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR3AHSX3_C_F_Z_R 0.1
`define NR3AHSX3_C_R_Z_F 0.1
`define NR3AHSX3_B_F_Z_R 0.1
`define NR3AHSX3_B_R_Z_F 0.1
`define NR3AHSX3_A_F_Z_F 0.1
`define NR3AHSX3_A_R_Z_R 0.1

module NR3AHSX3 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`NR3AHSX3_C_F_Z_R,`NR3AHSX3_C_R_Z_F);
      (B -=> Z) = (`NR3AHSX3_B_F_Z_R,`NR3AHSX3_B_R_Z_F);
      (A +=> Z) = (`NR3AHSX3_A_R_Z_R,`NR3AHSX3_A_F_Z_F);

   endspecify
`endif


endmodule // NR3AHSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:03 and Version :1.1 //
 
//  START 
// CELL NR3AHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR3AHSX4_C_F_Z_R 0.1
`define NR3AHSX4_C_R_Z_F 0.1
`define NR3AHSX4_B_F_Z_R 0.1
`define NR3AHSX4_B_R_Z_F 0.1
`define NR3AHSX4_A_F_Z_F 0.1
`define NR3AHSX4_A_R_Z_R 0.1

module NR3AHSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`NR3AHSX4_C_F_Z_R,`NR3AHSX4_C_R_Z_F);
      (B -=> Z) = (`NR3AHSX4_B_F_Z_R,`NR3AHSX4_B_R_Z_F);
      (A +=> Z) = (`NR3AHSX4_A_R_Z_R,`NR3AHSX4_A_F_Z_F);

   endspecify
`endif


endmodule // NR3AHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:03 and Version :1.1 //
 
//  START 
// CELL F_NR3AHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_NR3AHSP_C_F_Z_R 0.1
`define F_NR3AHSP_C_R_Z_F 0.1
`define F_NR3AHSP_B_F_Z_R 0.1
`define F_NR3AHSP_B_R_Z_F 0.1
`define F_NR3AHSP_A_F_Z_F 0.1
`define F_NR3AHSP_A_R_Z_R 0.1

module F_NR3AHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`F_NR3AHSP_C_F_Z_R,`F_NR3AHSP_C_R_Z_F);
      (B -=> Z) = (`F_NR3AHSP_B_F_Z_R,`F_NR3AHSP_B_R_Z_F);
      (A +=> Z) = (`F_NR3AHSP_A_R_Z_R,`F_NR3AHSP_A_F_Z_F);

   endspecify
`endif


endmodule // F_NR3AHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:03 and Version :1.1 //
 
//  START 
// CELL NR3AHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR3AHSX8_C_F_Z_R 0.1
`define NR3AHSX8_C_R_Z_F 0.1
`define NR3AHSX8_B_F_Z_R 0.1
`define NR3AHSX8_B_R_Z_F 0.1
`define NR3AHSX8_A_F_Z_F 0.1
`define NR3AHSX8_A_R_Z_R 0.1

module NR3AHSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   nor  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C -=> Z) = (`NR3AHSX8_C_F_Z_R,`NR3AHSX8_C_R_Z_F);
      (B -=> Z) = (`NR3AHSX8_B_F_Z_R,`NR3AHSX8_B_R_Z_F);
      (A +=> Z) = (`NR3AHSX8_A_R_Z_R,`NR3AHSX8_A_F_Z_F);

   endspecify
`endif


endmodule // NR3AHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:03 and Version :1.1 //
 
//  START 
// CELL NR4HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR4HSX05_D_F_Z_R 0.1
`define NR4HSX05_D_R_Z_F 0.1
`define NR4HSX05_C_F_Z_R 0.1
`define NR4HSX05_C_R_Z_F 0.1
`define NR4HSX05_B_F_Z_R 0.1
`define NR4HSX05_B_R_Z_F 0.1
`define NR4HSX05_A_F_Z_R 0.1
`define NR4HSX05_A_R_Z_F 0.1

module NR4HSX05 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`NR4HSX05_D_F_Z_R,`NR4HSX05_D_R_Z_F);
      (C -=> Z) = (`NR4HSX05_C_F_Z_R,`NR4HSX05_C_R_Z_F);
      (B -=> Z) = (`NR4HSX05_B_F_Z_R,`NR4HSX05_B_R_Z_F);
      (A -=> Z) = (`NR4HSX05_A_F_Z_R,`NR4HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // NR4HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:05 and Version :1.1 //
 
//  START 
// CELL NR4HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR4HS_D_F_Z_R 0.1
`define NR4HS_D_R_Z_F 0.1
`define NR4HS_C_F_Z_R 0.1
`define NR4HS_C_R_Z_F 0.1
`define NR4HS_B_F_Z_R 0.1
`define NR4HS_B_R_Z_F 0.1
`define NR4HS_A_F_Z_R 0.1
`define NR4HS_A_R_Z_F 0.1

module NR4HS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`NR4HS_D_F_Z_R,`NR4HS_D_R_Z_F);
      (C -=> Z) = (`NR4HS_C_F_Z_R,`NR4HS_C_R_Z_F);
      (B -=> Z) = (`NR4HS_B_F_Z_R,`NR4HS_B_R_Z_F);
      (A -=> Z) = (`NR4HS_A_F_Z_R,`NR4HS_A_R_Z_F);

   endspecify
`endif


endmodule // NR4HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:05 and Version :1.1 //
 
//  START 
// CELL NR4HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR4HSP_D_F_Z_R 0.1
`define NR4HSP_D_R_Z_F 0.1
`define NR4HSP_C_F_Z_R 0.1
`define NR4HSP_C_R_Z_F 0.1
`define NR4HSP_B_F_Z_R 0.1
`define NR4HSP_B_R_Z_F 0.1
`define NR4HSP_A_F_Z_R 0.1
`define NR4HSP_A_R_Z_F 0.1

module NR4HSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`NR4HSP_D_F_Z_R,`NR4HSP_D_R_Z_F);
      (C -=> Z) = (`NR4HSP_C_F_Z_R,`NR4HSP_C_R_Z_F);
      (B -=> Z) = (`NR4HSP_B_F_Z_R,`NR4HSP_B_R_Z_F);
      (A -=> Z) = (`NR4HSP_A_F_Z_R,`NR4HSP_A_R_Z_F);

   endspecify
`endif


endmodule // NR4HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:05 and Version :1.1 //
 
//  START 
// CELL NR4HSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR4HSX3_D_F_Z_R 0.1
`define NR4HSX3_D_R_Z_F 0.1
`define NR4HSX3_C_F_Z_R 0.1
`define NR4HSX3_C_R_Z_F 0.1
`define NR4HSX3_B_F_Z_R 0.1
`define NR4HSX3_B_R_Z_F 0.1
`define NR4HSX3_A_F_Z_R 0.1
`define NR4HSX3_A_R_Z_F 0.1

module NR4HSX3 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`NR4HSX3_D_F_Z_R,`NR4HSX3_D_R_Z_F);
      (C -=> Z) = (`NR4HSX3_C_F_Z_R,`NR4HSX3_C_R_Z_F);
      (B -=> Z) = (`NR4HSX3_B_F_Z_R,`NR4HSX3_B_R_Z_F);
      (A -=> Z) = (`NR4HSX3_A_F_Z_R,`NR4HSX3_A_R_Z_F);

   endspecify
`endif


endmodule // NR4HSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:05 and Version :1.1 //
 
//  START 
// CELL NR4HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR4HSX4_D_F_Z_R 0.1
`define NR4HSX4_D_R_Z_F 0.1
`define NR4HSX4_C_F_Z_R 0.1
`define NR4HSX4_C_R_Z_F 0.1
`define NR4HSX4_B_F_Z_R 0.1
`define NR4HSX4_B_R_Z_F 0.1
`define NR4HSX4_A_F_Z_R 0.1
`define NR4HSX4_A_R_Z_F 0.1

module NR4HSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`NR4HSX4_D_F_Z_R,`NR4HSX4_D_R_Z_F);
      (C -=> Z) = (`NR4HSX4_C_F_Z_R,`NR4HSX4_C_R_Z_F);
      (B -=> Z) = (`NR4HSX4_B_F_Z_R,`NR4HSX4_B_R_Z_F);
      (A -=> Z) = (`NR4HSX4_A_F_Z_R,`NR4HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // NR4HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:05 and Version :1.1 //
 
//  START 
// CELL NR4HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR4HSX8_D_F_Z_R 0.1
`define NR4HSX8_D_R_Z_F 0.1
`define NR4HSX8_C_F_Z_R 0.1
`define NR4HSX8_C_R_Z_F 0.1
`define NR4HSX8_B_F_Z_R 0.1
`define NR4HSX8_B_R_Z_F 0.1
`define NR4HSX8_A_F_Z_R 0.1
`define NR4HSX8_A_R_Z_F 0.1

module NR4HSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`NR4HSX8_D_F_Z_R,`NR4HSX8_D_R_Z_F);
      (C -=> Z) = (`NR4HSX8_C_F_Z_R,`NR4HSX8_C_R_Z_F);
      (B -=> Z) = (`NR4HSX8_B_F_Z_R,`NR4HSX8_B_R_Z_F);
      (A -=> Z) = (`NR4HSX8_A_F_Z_R,`NR4HSX8_A_R_Z_F);

   endspecify
`endif


endmodule // NR4HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:05 and Version :1.1 //
 
//  START 
// CELL F_NR4HSX05

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_NR4HSX05_D_F_Z_R 0.1
`define F_NR4HSX05_D_R_Z_F 0.1
`define F_NR4HSX05_C_F_Z_R 0.1
`define F_NR4HSX05_C_R_Z_F 0.1
`define F_NR4HSX05_B_F_Z_R 0.1
`define F_NR4HSX05_B_R_Z_F 0.1
`define F_NR4HSX05_A_F_Z_R 0.1
`define F_NR4HSX05_A_R_Z_F 0.1

module F_NR4HSX05 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   nor  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D -=> Z) = (`F_NR4HSX05_D_F_Z_R,`F_NR4HSX05_D_R_Z_F);
      (C -=> Z) = (`F_NR4HSX05_C_F_Z_R,`F_NR4HSX05_C_R_Z_F);
      (B -=> Z) = (`F_NR4HSX05_B_F_Z_R,`F_NR4HSX05_B_R_Z_F);
      (A -=> Z) = (`F_NR4HSX05_A_F_Z_R,`F_NR4HSX05_A_R_Z_F);

   endspecify
`endif


endmodule // F_NR4HSX05
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:05 and Version :1.1 //
 
//  START 
// CELL NR5HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR5HS_E_F_Z_R 0.1
`define NR5HS_E_R_Z_F 0.1
`define NR5HS_D_F_Z_R 0.1
`define NR5HS_D_R_Z_F 0.1
`define NR5HS_C_F_Z_R 0.1
`define NR5HS_C_R_Z_F 0.1
`define NR5HS_B_F_Z_R 0.1
`define NR5HS_B_R_Z_F 0.1
`define NR5HS_A_F_Z_R 0.1
`define NR5HS_A_R_Z_F 0.1

module NR5HS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   nor  u0 (Z, A, B, C, D, E);


`ifdef functional
`else
   specify

      (E -=> Z) = (`NR5HS_E_F_Z_R,`NR5HS_E_R_Z_F);
      (D -=> Z) = (`NR5HS_D_F_Z_R,`NR5HS_D_R_Z_F);
      (C -=> Z) = (`NR5HS_C_F_Z_R,`NR5HS_C_R_Z_F);
      (B -=> Z) = (`NR5HS_B_F_Z_R,`NR5HS_B_R_Z_F);
      (A -=> Z) = (`NR5HS_A_F_Z_R,`NR5HS_A_R_Z_F);

   endspecify
`endif


endmodule // NR5HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:11 and Version :1.1 //
 
//  START 
// CELL NR5HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR5HSP_E_F_Z_R 0.1
`define NR5HSP_E_R_Z_F 0.1
`define NR5HSP_D_F_Z_R 0.1
`define NR5HSP_D_R_Z_F 0.1
`define NR5HSP_C_F_Z_R 0.1
`define NR5HSP_C_R_Z_F 0.1
`define NR5HSP_B_F_Z_R 0.1
`define NR5HSP_B_R_Z_F 0.1
`define NR5HSP_A_F_Z_R 0.1
`define NR5HSP_A_R_Z_F 0.1

module NR5HSP (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   nor  u0 (Z, A, B, C, D, E);


`ifdef functional
`else
   specify

      (E -=> Z) = (`NR5HSP_E_F_Z_R,`NR5HSP_E_R_Z_F);
      (D -=> Z) = (`NR5HSP_D_F_Z_R,`NR5HSP_D_R_Z_F);
      (C -=> Z) = (`NR5HSP_C_F_Z_R,`NR5HSP_C_R_Z_F);
      (B -=> Z) = (`NR5HSP_B_F_Z_R,`NR5HSP_B_R_Z_F);
      (A -=> Z) = (`NR5HSP_A_F_Z_R,`NR5HSP_A_R_Z_F);

   endspecify
`endif


endmodule // NR5HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:11 and Version :1.1 //
 
//  START 
// CELL NR5HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR5HSX4_E_F_Z_R 0.1
`define NR5HSX4_E_R_Z_F 0.1
`define NR5HSX4_D_F_Z_R 0.1
`define NR5HSX4_D_R_Z_F 0.1
`define NR5HSX4_C_F_Z_R 0.1
`define NR5HSX4_C_R_Z_F 0.1
`define NR5HSX4_B_F_Z_R 0.1
`define NR5HSX4_B_R_Z_F 0.1
`define NR5HSX4_A_F_Z_R 0.1
`define NR5HSX4_A_R_Z_F 0.1

module NR5HSX4 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   nor  u0 (Z, A, B, C, D, E);


`ifdef functional
`else
   specify

      (E -=> Z) = (`NR5HSX4_E_F_Z_R,`NR5HSX4_E_R_Z_F);
      (D -=> Z) = (`NR5HSX4_D_F_Z_R,`NR5HSX4_D_R_Z_F);
      (C -=> Z) = (`NR5HSX4_C_F_Z_R,`NR5HSX4_C_R_Z_F);
      (B -=> Z) = (`NR5HSX4_B_F_Z_R,`NR5HSX4_B_R_Z_F);
      (A -=> Z) = (`NR5HSX4_A_F_Z_R,`NR5HSX4_A_R_Z_F);

   endspecify
`endif


endmodule // NR5HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:11 and Version :1.1 //
 
//  START 
// CELL NR6HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR6HS_F_F_Z_R 0.1
`define NR6HS_F_R_Z_F 0.1
`define NR6HS_E_F_Z_R 0.1
`define NR6HS_E_R_Z_F 0.1
`define NR6HS_D_F_Z_R 0.1
`define NR6HS_D_R_Z_F 0.1
`define NR6HS_C_F_Z_R 0.1
`define NR6HS_C_R_Z_F 0.1
`define NR6HS_B_F_Z_R 0.1
`define NR6HS_B_R_Z_F 0.1
`define NR6HS_A_F_Z_R 0.1
`define NR6HS_A_R_Z_F 0.1

module NR6HS (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   nor  u0 (Z, A, B, C, D, E, F);


`ifdef functional
`else
   specify

      (F -=> Z) = (`NR6HS_F_F_Z_R,`NR6HS_F_R_Z_F);
      (E -=> Z) = (`NR6HS_E_F_Z_R,`NR6HS_E_R_Z_F);
      (D -=> Z) = (`NR6HS_D_F_Z_R,`NR6HS_D_R_Z_F);
      (C -=> Z) = (`NR6HS_C_F_Z_R,`NR6HS_C_R_Z_F);
      (B -=> Z) = (`NR6HS_B_F_Z_R,`NR6HS_B_R_Z_F);
      (A -=> Z) = (`NR6HS_A_F_Z_R,`NR6HS_A_R_Z_F);

   endspecify
`endif


endmodule // NR6HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:18 and Version :1.1 //
 
//  START 
// CELL NR7HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR7HS_G_F_Z_R 0.1
`define NR7HS_G_R_Z_F 0.1
`define NR7HS_F_F_Z_R 0.1
`define NR7HS_F_R_Z_F 0.1
`define NR7HS_E_F_Z_R 0.1
`define NR7HS_E_R_Z_F 0.1
`define NR7HS_D_F_Z_R 0.1
`define NR7HS_D_R_Z_F 0.1
`define NR7HS_C_F_Z_R 0.1
`define NR7HS_C_R_Z_F 0.1
`define NR7HS_B_F_Z_R 0.1
`define NR7HS_B_R_Z_F 0.1
`define NR7HS_A_F_Z_R 0.1
`define NR7HS_A_R_Z_F 0.1

module NR7HS (Z, A, B, C, D, E, F, G);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;
   input G;


   nor  u0 (Z, A, B, C, D, E, F, G);


`ifdef functional
`else
   specify

      (G -=> Z) = (`NR7HS_G_F_Z_R,`NR7HS_G_R_Z_F);
      (F -=> Z) = (`NR7HS_F_F_Z_R,`NR7HS_F_R_Z_F);
      (E -=> Z) = (`NR7HS_E_F_Z_R,`NR7HS_E_R_Z_F);
      (D -=> Z) = (`NR7HS_D_F_Z_R,`NR7HS_D_R_Z_F);
      (C -=> Z) = (`NR7HS_C_F_Z_R,`NR7HS_C_R_Z_F);
      (B -=> Z) = (`NR7HS_B_F_Z_R,`NR7HS_B_R_Z_F);
      (A -=> Z) = (`NR7HS_A_F_Z_R,`NR7HS_A_R_Z_F);

   endspecify
`endif


endmodule // NR7HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:22 and Version :1.1 //
 
//  START 
// CELL NR8HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define NR8HS_H_F_Z_R 0.1
`define NR8HS_H_R_Z_F 0.1
`define NR8HS_G_F_Z_R 0.1
`define NR8HS_G_R_Z_F 0.1
`define NR8HS_F_F_Z_R 0.1
`define NR8HS_F_R_Z_F 0.1
`define NR8HS_E_F_Z_R 0.1
`define NR8HS_E_R_Z_F 0.1
`define NR8HS_D_F_Z_R 0.1
`define NR8HS_D_R_Z_F 0.1
`define NR8HS_C_F_Z_R 0.1
`define NR8HS_C_R_Z_F 0.1
`define NR8HS_B_F_Z_R 0.1
`define NR8HS_B_R_Z_F 0.1
`define NR8HS_A_F_Z_R 0.1
`define NR8HS_A_R_Z_F 0.1

module NR8HS (Z, A, B, C, D, E, F, G, H);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;
   input G;
   input H;


   nor  u0 (Z, A, B, C, D, E, F, G, H);


`ifdef functional
`else
   specify

      (H -=> Z) = (`NR8HS_H_F_Z_R,`NR8HS_H_R_Z_F);
      (G -=> Z) = (`NR8HS_G_F_Z_R,`NR8HS_G_R_Z_F);
      (F -=> Z) = (`NR8HS_F_F_Z_R,`NR8HS_F_R_Z_F);
      (E -=> Z) = (`NR8HS_E_F_Z_R,`NR8HS_E_R_Z_F);
      (D -=> Z) = (`NR8HS_D_F_Z_R,`NR8HS_D_R_Z_F);
      (C -=> Z) = (`NR8HS_C_F_Z_R,`NR8HS_C_R_Z_F);
      (B -=> Z) = (`NR8HS_B_F_Z_R,`NR8HS_B_R_Z_F);
      (A -=> Z) = (`NR8HS_A_F_Z_R,`NR8HS_A_R_Z_F);

   endspecify
`endif


endmodule // NR8HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:25 and Version :1.1 //
 
//  START 
// CELL OR2HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR2HS_B_F_Z_F 0.1
`define OR2HS_B_R_Z_R 0.1
`define OR2HS_A_F_Z_F 0.1
`define OR2HS_A_R_Z_R 0.1

module OR2HS (Z, A, B);

   output Z;
   input A;
   input B;


   or  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B +=> Z) = (`OR2HS_B_R_Z_R,`OR2HS_B_F_Z_F);
      (A +=> Z) = (`OR2HS_A_R_Z_R,`OR2HS_A_F_Z_F);

   endspecify
`endif


endmodule // OR2HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:27 and Version :1.1 //
 
//  START 
// CELL OR2HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR2HSP_B_F_Z_F 0.1
`define OR2HSP_B_R_Z_R 0.1
`define OR2HSP_A_F_Z_F 0.1
`define OR2HSP_A_R_Z_R 0.1

module OR2HSP (Z, A, B);

   output Z;
   input A;
   input B;


   or  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B +=> Z) = (`OR2HSP_B_R_Z_R,`OR2HSP_B_F_Z_F);
      (A +=> Z) = (`OR2HSP_A_R_Z_R,`OR2HSP_A_F_Z_F);

   endspecify
`endif


endmodule // OR2HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:27 and Version :1.1 //
 
//  START 
// CELL OR2HSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR2HSX3_B_F_Z_F 0.1
`define OR2HSX3_B_R_Z_R 0.1
`define OR2HSX3_A_F_Z_F 0.1
`define OR2HSX3_A_R_Z_R 0.1

module OR2HSX3 (Z, A, B);

   output Z;
   input A;
   input B;


   or  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B +=> Z) = (`OR2HSX3_B_R_Z_R,`OR2HSX3_B_F_Z_F);
      (A +=> Z) = (`OR2HSX3_A_R_Z_R,`OR2HSX3_A_F_Z_F);

   endspecify
`endif


endmodule // OR2HSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:27 and Version :1.1 //
 
//  START 
// CELL OR2HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR2HSX4_B_F_Z_F 0.1
`define OR2HSX4_B_R_Z_R 0.1
`define OR2HSX4_A_F_Z_F 0.1
`define OR2HSX4_A_R_Z_R 0.1

module OR2HSX4 (Z, A, B);

   output Z;
   input A;
   input B;


   or  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B +=> Z) = (`OR2HSX4_B_R_Z_R,`OR2HSX4_B_F_Z_F);
      (A +=> Z) = (`OR2HSX4_A_R_Z_R,`OR2HSX4_A_F_Z_F);

   endspecify
`endif


endmodule // OR2HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:27 and Version :1.1 //
 
//  START 
// CELL OR2HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR2HSX8_B_F_Z_F 0.1
`define OR2HSX8_B_R_Z_R 0.1
`define OR2HSX8_A_F_Z_F 0.1
`define OR2HSX8_A_R_Z_R 0.1

module OR2HSX8 (Z, A, B);

   output Z;
   input A;
   input B;


   or  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B +=> Z) = (`OR2HSX8_B_R_Z_R,`OR2HSX8_B_F_Z_F);
      (A +=> Z) = (`OR2HSX8_A_R_Z_R,`OR2HSX8_A_F_Z_F);

   endspecify
`endif


endmodule // OR2HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:27 and Version :1.1 //
 
//  START 
// CELL F_OR2HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_OR2HSX4_B_F_Z_F 0.1
`define F_OR2HSX4_B_R_Z_R 0.1
`define F_OR2HSX4_A_F_Z_F 0.1
`define F_OR2HSX4_A_R_Z_R 0.1

module F_OR2HSX4 (Z, A, B);

   output Z;
   input A;
   input B;


   or  u0 (Z, A, B);


`ifdef functional
`else
   specify

      (B +=> Z) = (`F_OR2HSX4_B_R_Z_R,`F_OR2HSX4_B_F_Z_F);
      (A +=> Z) = (`F_OR2HSX4_A_R_Z_R,`F_OR2HSX4_A_F_Z_F);

   endspecify
`endif


endmodule // F_OR2HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:27 and Version :1.1 //
 
//  START 
// CELL OR2AHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR2AHS_B_F_Z_F 0.1
`define OR2AHS_B_R_Z_R 0.1
`define OR2AHS_A_F_Z_R 0.1
`define OR2AHS_A_R_Z_F 0.1

module OR2AHS (Z, A, B);

   output Z;
   input A;
   input B;


   or  u0 (Z, AX, B);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (B +=> Z) = (`OR2AHS_B_R_Z_R,`OR2AHS_B_F_Z_F);
      (A -=> Z) = (`OR2AHS_A_F_Z_R,`OR2AHS_A_R_Z_F);

   endspecify
`endif


endmodule // OR2AHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:27 and Version :1.1 //
 
//  START 
// CELL OR2AHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR2AHSP_B_F_Z_F 0.1
`define OR2AHSP_B_R_Z_R 0.1
`define OR2AHSP_A_F_Z_R 0.1
`define OR2AHSP_A_R_Z_F 0.1

module OR2AHSP (Z, A, B);

   output Z;
   input A;
   input B;


   or  u0 (Z, AX, B);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (B +=> Z) = (`OR2AHSP_B_R_Z_R,`OR2AHSP_B_F_Z_F);
      (A -=> Z) = (`OR2AHSP_A_F_Z_R,`OR2AHSP_A_R_Z_F);

   endspecify
`endif


endmodule // OR2AHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:27 and Version :1.1 //
 
//  START 
// CELL OR2AHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR2AHSX4_B_F_Z_F 0.1
`define OR2AHSX4_B_R_Z_R 0.1
`define OR2AHSX4_A_F_Z_R 0.1
`define OR2AHSX4_A_R_Z_F 0.1

module OR2AHSX4 (Z, A, B);

   output Z;
   input A;
   input B;


   or  u0 (Z, AX, B);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (B +=> Z) = (`OR2AHSX4_B_R_Z_R,`OR2AHSX4_B_F_Z_F);
      (A -=> Z) = (`OR2AHSX4_A_F_Z_R,`OR2AHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // OR2AHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:27 and Version :1.1 //
 
//  START 
// CELL OR2AHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR2AHSX8_B_F_Z_F 0.1
`define OR2AHSX8_B_R_Z_R 0.1
`define OR2AHSX8_A_F_Z_R 0.1
`define OR2AHSX8_A_R_Z_F 0.1

module OR2AHSX8 (Z, A, B);

   output Z;
   input A;
   input B;


   or  u0 (Z, AX, B);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (B +=> Z) = (`OR2AHSX8_B_R_Z_R,`OR2AHSX8_B_F_Z_F);
      (A -=> Z) = (`OR2AHSX8_A_F_Z_R,`OR2AHSX8_A_R_Z_F);

   endspecify
`endif


endmodule // OR2AHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:27 and Version :1.1 //
 
//  START 
// CELL OR3HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR3HS_C_F_Z_F 0.1
`define OR3HS_C_R_Z_R 0.1
`define OR3HS_B_F_Z_F 0.1
`define OR3HS_B_R_Z_R 0.1
`define OR3HS_A_F_Z_F 0.1
`define OR3HS_A_R_Z_R 0.1

module OR3HS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C +=> Z) = (`OR3HS_C_R_Z_R,`OR3HS_C_F_Z_F);
      (B +=> Z) = (`OR3HS_B_R_Z_R,`OR3HS_B_F_Z_F);
      (A +=> Z) = (`OR3HS_A_R_Z_R,`OR3HS_A_F_Z_F);

   endspecify
`endif


endmodule // OR3HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:33 and Version :1.1 //
 
//  START 
// CELL OR3HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR3HSP_C_F_Z_F 0.1
`define OR3HSP_C_R_Z_R 0.1
`define OR3HSP_B_F_Z_F 0.1
`define OR3HSP_B_R_Z_R 0.1
`define OR3HSP_A_F_Z_F 0.1
`define OR3HSP_A_R_Z_R 0.1

module OR3HSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C +=> Z) = (`OR3HSP_C_R_Z_R,`OR3HSP_C_F_Z_F);
      (B +=> Z) = (`OR3HSP_B_R_Z_R,`OR3HSP_B_F_Z_F);
      (A +=> Z) = (`OR3HSP_A_R_Z_R,`OR3HSP_A_F_Z_F);

   endspecify
`endif


endmodule // OR3HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:33 and Version :1.1 //
 
//  START 
// CELL OR3HSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR3HSX3_C_F_Z_F 0.1
`define OR3HSX3_C_R_Z_R 0.1
`define OR3HSX3_B_F_Z_F 0.1
`define OR3HSX3_B_R_Z_R 0.1
`define OR3HSX3_A_F_Z_F 0.1
`define OR3HSX3_A_R_Z_R 0.1

module OR3HSX3 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C +=> Z) = (`OR3HSX3_C_R_Z_R,`OR3HSX3_C_F_Z_F);
      (B +=> Z) = (`OR3HSX3_B_R_Z_R,`OR3HSX3_B_F_Z_F);
      (A +=> Z) = (`OR3HSX3_A_R_Z_R,`OR3HSX3_A_F_Z_F);

   endspecify
`endif


endmodule // OR3HSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:33 and Version :1.1 //
 
//  START 
// CELL OR3HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR3HSX4_C_F_Z_F 0.1
`define OR3HSX4_C_R_Z_R 0.1
`define OR3HSX4_B_F_Z_F 0.1
`define OR3HSX4_B_R_Z_R 0.1
`define OR3HSX4_A_F_Z_F 0.1
`define OR3HSX4_A_R_Z_R 0.1

module OR3HSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C +=> Z) = (`OR3HSX4_C_R_Z_R,`OR3HSX4_C_F_Z_F);
      (B +=> Z) = (`OR3HSX4_B_R_Z_R,`OR3HSX4_B_F_Z_F);
      (A +=> Z) = (`OR3HSX4_A_R_Z_R,`OR3HSX4_A_F_Z_F);

   endspecify
`endif


endmodule // OR3HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:33 and Version :1.1 //
 
//  START 
// CELL F_OR3HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define F_OR3HSX4_C_F_Z_F 0.1
`define F_OR3HSX4_C_R_Z_R 0.1
`define F_OR3HSX4_B_F_Z_F 0.1
`define F_OR3HSX4_B_R_Z_R 0.1
`define F_OR3HSX4_A_F_Z_F 0.1
`define F_OR3HSX4_A_R_Z_R 0.1

module F_OR3HSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C +=> Z) = (`F_OR3HSX4_C_R_Z_R,`F_OR3HSX4_C_F_Z_F);
      (B +=> Z) = (`F_OR3HSX4_B_R_Z_R,`F_OR3HSX4_B_F_Z_F);
      (A +=> Z) = (`F_OR3HSX4_A_R_Z_R,`F_OR3HSX4_A_F_Z_F);

   endspecify
`endif


endmodule // F_OR3HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:33 and Version :1.1 //
 
//  START 
// CELL OR3HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR3HSX8_C_F_Z_F 0.1
`define OR3HSX8_C_R_Z_R 0.1
`define OR3HSX8_B_F_Z_F 0.1
`define OR3HSX8_B_R_Z_R 0.1
`define OR3HSX8_A_F_Z_F 0.1
`define OR3HSX8_A_R_Z_R 0.1

module OR3HSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, A, B, C);


`ifdef functional
`else
   specify

      (C +=> Z) = (`OR3HSX8_C_R_Z_R,`OR3HSX8_C_F_Z_F);
      (B +=> Z) = (`OR3HSX8_B_R_Z_R,`OR3HSX8_B_F_Z_F);
      (A +=> Z) = (`OR3HSX8_A_R_Z_R,`OR3HSX8_A_F_Z_F);

   endspecify
`endif


endmodule // OR3HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:33 and Version :1.1 //
 
//  START 
// CELL OR3AHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR3AHS_C_F_Z_F 0.1
`define OR3AHS_C_R_Z_R 0.1
`define OR3AHS_B_F_Z_F 0.1
`define OR3AHS_B_R_Z_R 0.1
`define OR3AHS_A_F_Z_R 0.1
`define OR3AHS_A_R_Z_F 0.1

module OR3AHS (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C +=> Z) = (`OR3AHS_C_R_Z_R,`OR3AHS_C_F_Z_F);
      (B +=> Z) = (`OR3AHS_B_R_Z_R,`OR3AHS_B_F_Z_F);
      (A -=> Z) = (`OR3AHS_A_F_Z_R,`OR3AHS_A_R_Z_F);

   endspecify
`endif


endmodule // OR3AHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:33 and Version :1.1 //
 
//  START 
// CELL OR3AHSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR3AHSP_C_F_Z_F 0.1
`define OR3AHSP_C_R_Z_R 0.1
`define OR3AHSP_B_F_Z_F 0.1
`define OR3AHSP_B_R_Z_R 0.1
`define OR3AHSP_A_F_Z_R 0.1
`define OR3AHSP_A_R_Z_F 0.1

module OR3AHSP (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C +=> Z) = (`OR3AHSP_C_R_Z_R,`OR3AHSP_C_F_Z_F);
      (B +=> Z) = (`OR3AHSP_B_R_Z_R,`OR3AHSP_B_F_Z_F);
      (A -=> Z) = (`OR3AHSP_A_F_Z_R,`OR3AHSP_A_R_Z_F);

   endspecify
`endif


endmodule // OR3AHSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:33 and Version :1.1 //
 
//  START 
// CELL OR3AHSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR3AHSX3_C_F_Z_F 0.1
`define OR3AHSX3_C_R_Z_R 0.1
`define OR3AHSX3_B_F_Z_F 0.1
`define OR3AHSX3_B_R_Z_R 0.1
`define OR3AHSX3_A_F_Z_R 0.1
`define OR3AHSX3_A_R_Z_F 0.1

module OR3AHSX3 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C +=> Z) = (`OR3AHSX3_C_R_Z_R,`OR3AHSX3_C_F_Z_F);
      (B +=> Z) = (`OR3AHSX3_B_R_Z_R,`OR3AHSX3_B_F_Z_F);
      (A -=> Z) = (`OR3AHSX3_A_F_Z_R,`OR3AHSX3_A_R_Z_F);

   endspecify
`endif


endmodule // OR3AHSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:33 and Version :1.1 //
 
//  START 
// CELL OR3AHSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR3AHSX4_C_F_Z_F 0.1
`define OR3AHSX4_C_R_Z_R 0.1
`define OR3AHSX4_B_F_Z_F 0.1
`define OR3AHSX4_B_R_Z_R 0.1
`define OR3AHSX4_A_F_Z_R 0.1
`define OR3AHSX4_A_R_Z_F 0.1

module OR3AHSX4 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C +=> Z) = (`OR3AHSX4_C_R_Z_R,`OR3AHSX4_C_F_Z_F);
      (B +=> Z) = (`OR3AHSX4_B_R_Z_R,`OR3AHSX4_B_F_Z_F);
      (A -=> Z) = (`OR3AHSX4_A_F_Z_R,`OR3AHSX4_A_R_Z_F);

   endspecify
`endif


endmodule // OR3AHSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:33 and Version :1.1 //
 
//  START 
// CELL OR3AHSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR3AHSX8_C_F_Z_F 0.1
`define OR3AHSX8_C_R_Z_R 0.1
`define OR3AHSX8_B_F_Z_F 0.1
`define OR3AHSX8_B_R_Z_R 0.1
`define OR3AHSX8_A_F_Z_R 0.1
`define OR3AHSX8_A_R_Z_F 0.1

module OR3AHSX8 (Z, A, B, C);

   output Z;
   input A;
   input B;
   input C;


   or  u0 (Z, AX, B, C);
   not  u1 (AX, A);


`ifdef functional
`else
   specify

      (C +=> Z) = (`OR3AHSX8_C_R_Z_R,`OR3AHSX8_C_F_Z_F);
      (B +=> Z) = (`OR3AHSX8_B_R_Z_R,`OR3AHSX8_B_F_Z_F);
      (A -=> Z) = (`OR3AHSX8_A_F_Z_R,`OR3AHSX8_A_R_Z_F);

   endspecify
`endif


endmodule // OR3AHSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:33 and Version :1.1 //
 
//  START 
// CELL OR4HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR4HS_D_F_Z_F 0.1
`define OR4HS_D_R_Z_R 0.1
`define OR4HS_C_F_Z_F 0.1
`define OR4HS_C_R_Z_R 0.1
`define OR4HS_B_F_Z_F 0.1
`define OR4HS_B_R_Z_R 0.1
`define OR4HS_A_F_Z_F 0.1
`define OR4HS_A_R_Z_R 0.1

module OR4HS (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`OR4HS_D_R_Z_R,`OR4HS_D_F_Z_F);
      (C +=> Z) = (`OR4HS_C_R_Z_R,`OR4HS_C_F_Z_F);
      (B +=> Z) = (`OR4HS_B_R_Z_R,`OR4HS_B_F_Z_F);
      (A +=> Z) = (`OR4HS_A_R_Z_R,`OR4HS_A_F_Z_F);

   endspecify
`endif


endmodule // OR4HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:37 and Version :1.1 //
 
 
//  START
 


// CELL OR4HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR4HSP_D_F_Z_F 0.1
`define OR4HSP_D_R_Z_R 0.1
`define OR4HSP_C_F_Z_F 0.1
`define OR4HSP_C_R_Z_R 0.1
`define OR4HSP_B_F_Z_F 0.1
`define OR4HSP_B_R_Z_R 0.1
`define OR4HSP_A_F_Z_F 0.1
`define OR4HSP_A_R_Z_R 0.1

module OR4HSP (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`OR4HSP_D_R_Z_R,`OR4HSP_D_F_Z_F);
      (C +=> Z) = (`OR4HSP_C_R_Z_R,`OR4HSP_C_F_Z_F);
      (B +=> Z) = (`OR4HSP_B_R_Z_R,`OR4HSP_B_F_Z_F);
      (A +=> Z) = (`OR4HSP_A_R_Z_R,`OR4HSP_A_F_Z_F);

   endspecify
`endif


endmodule // OR4HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:37 and Version :1.1 //
 
 
//  START
 


// CELL OR4HSX3

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR4HSX3_D_F_Z_F 0.1
`define OR4HSX3_D_R_Z_R 0.1
`define OR4HSX3_C_F_Z_F 0.1
`define OR4HSX3_C_R_Z_R 0.1
`define OR4HSX3_B_F_Z_F 0.1
`define OR4HSX3_B_R_Z_R 0.1
`define OR4HSX3_A_F_Z_F 0.1
`define OR4HSX3_A_R_Z_R 0.1

module OR4HSX3 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`OR4HSX3_D_R_Z_R,`OR4HSX3_D_F_Z_F);
      (C +=> Z) = (`OR4HSX3_C_R_Z_R,`OR4HSX3_C_F_Z_F);
      (B +=> Z) = (`OR4HSX3_B_R_Z_R,`OR4HSX3_B_F_Z_F);
      (A +=> Z) = (`OR4HSX3_A_R_Z_R,`OR4HSX3_A_F_Z_F);

   endspecify
`endif


endmodule // OR4HSX3
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:37 and Version :1.1 //
 
 
//  START
 


// CELL OR4HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR4HSX4_D_F_Z_F 0.1
`define OR4HSX4_D_R_Z_R 0.1
`define OR4HSX4_C_F_Z_F 0.1
`define OR4HSX4_C_R_Z_R 0.1
`define OR4HSX4_B_F_Z_F 0.1
`define OR4HSX4_B_R_Z_R 0.1
`define OR4HSX4_A_F_Z_F 0.1
`define OR4HSX4_A_R_Z_R 0.1

module OR4HSX4 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`OR4HSX4_D_R_Z_R,`OR4HSX4_D_F_Z_F);
      (C +=> Z) = (`OR4HSX4_C_R_Z_R,`OR4HSX4_C_F_Z_F);
      (B +=> Z) = (`OR4HSX4_B_R_Z_R,`OR4HSX4_B_F_Z_F);
      (A +=> Z) = (`OR4HSX4_A_R_Z_R,`OR4HSX4_A_F_Z_F);

   endspecify
`endif


endmodule // OR4HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:37 and Version :1.1 //
 
 
//  START
 


// CELL OR4HSX8

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR4HSX8_D_F_Z_F 0.1
`define OR4HSX8_D_R_Z_R 0.1
`define OR4HSX8_C_F_Z_F 0.1
`define OR4HSX8_C_R_Z_R 0.1
`define OR4HSX8_B_F_Z_F 0.1
`define OR4HSX8_B_R_Z_R 0.1
`define OR4HSX8_A_F_Z_F 0.1
`define OR4HSX8_A_R_Z_R 0.1

module OR4HSX8 (Z, A, B, C, D);

   output Z;
   input A;
   input B;
   input C;
   input D;


   or  u0 (Z, A, B, C, D);


`ifdef functional
`else
   specify

      (D +=> Z) = (`OR4HSX8_D_R_Z_R,`OR4HSX8_D_F_Z_F);
      (C +=> Z) = (`OR4HSX8_C_R_Z_R,`OR4HSX8_C_F_Z_F);
      (B +=> Z) = (`OR4HSX8_B_R_Z_R,`OR4HSX8_B_F_Z_F);
      (A +=> Z) = (`OR4HSX8_A_R_Z_R,`OR4HSX8_A_F_Z_F);

   endspecify
`endif


endmodule // OR4HSX8
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:37 and Version :1.1 //
 
 
//  START
 


// CELL OR5HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR5HS_E_F_Z_F 0.1
`define OR5HS_E_R_Z_R 0.1
`define OR5HS_D_F_Z_F 0.1
`define OR5HS_D_R_Z_R 0.1
`define OR5HS_C_F_Z_F 0.1
`define OR5HS_C_R_Z_R 0.1
`define OR5HS_B_F_Z_F 0.1
`define OR5HS_B_R_Z_R 0.1
`define OR5HS_A_F_Z_F 0.1
`define OR5HS_A_R_Z_R 0.1

module OR5HS (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   or  u0 (Z, A, B, C, D, E);


`ifdef functional
`else
   specify

      (E +=> Z) = (`OR5HS_E_R_Z_R,`OR5HS_E_F_Z_F);
      (D +=> Z) = (`OR5HS_D_R_Z_R,`OR5HS_D_F_Z_F);
      (C +=> Z) = (`OR5HS_C_R_Z_R,`OR5HS_C_F_Z_F);
      (B +=> Z) = (`OR5HS_B_R_Z_R,`OR5HS_B_F_Z_F);
      (A +=> Z) = (`OR5HS_A_R_Z_R,`OR5HS_A_F_Z_F);

   endspecify
`endif


endmodule // OR5HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:44 and Version :1.1 //
 
//  START 
// CELL OR5HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR5HSP_E_F_Z_F 0.1
`define OR5HSP_E_R_Z_R 0.1
`define OR5HSP_D_F_Z_F 0.1
`define OR5HSP_D_R_Z_R 0.1
`define OR5HSP_C_F_Z_F 0.1
`define OR5HSP_C_R_Z_R 0.1
`define OR5HSP_B_F_Z_F 0.1
`define OR5HSP_B_R_Z_R 0.1
`define OR5HSP_A_F_Z_F 0.1
`define OR5HSP_A_R_Z_R 0.1

module OR5HSP (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   or  u0 (Z, A, B, C, D, E);


`ifdef functional
`else
   specify

      (E +=> Z) = (`OR5HSP_E_R_Z_R,`OR5HSP_E_F_Z_F);
      (D +=> Z) = (`OR5HSP_D_R_Z_R,`OR5HSP_D_F_Z_F);
      (C +=> Z) = (`OR5HSP_C_R_Z_R,`OR5HSP_C_F_Z_F);
      (B +=> Z) = (`OR5HSP_B_R_Z_R,`OR5HSP_B_F_Z_F);
      (A +=> Z) = (`OR5HSP_A_R_Z_R,`OR5HSP_A_F_Z_F);

   endspecify
`endif


endmodule // OR5HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:44 and Version :1.1 //
 
//  START 
// CELL OR5HSX4

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR5HSX4_E_F_Z_F 0.1
`define OR5HSX4_E_R_Z_R 0.1
`define OR5HSX4_D_F_Z_F 0.1
`define OR5HSX4_D_R_Z_R 0.1
`define OR5HSX4_C_F_Z_F 0.1
`define OR5HSX4_C_R_Z_R 0.1
`define OR5HSX4_B_F_Z_F 0.1
`define OR5HSX4_B_R_Z_R 0.1
`define OR5HSX4_A_F_Z_F 0.1
`define OR5HSX4_A_R_Z_R 0.1

module OR5HSX4 (Z, A, B, C, D, E);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;


   or  u0 (Z, A, B, C, D, E);


`ifdef functional
`else
   specify

      (E +=> Z) = (`OR5HSX4_E_R_Z_R,`OR5HSX4_E_F_Z_F);
      (D +=> Z) = (`OR5HSX4_D_R_Z_R,`OR5HSX4_D_F_Z_F);
      (C +=> Z) = (`OR5HSX4_C_R_Z_R,`OR5HSX4_C_F_Z_F);
      (B +=> Z) = (`OR5HSX4_B_R_Z_R,`OR5HSX4_B_F_Z_F);
      (A +=> Z) = (`OR5HSX4_A_R_Z_R,`OR5HSX4_A_F_Z_F);

   endspecify
`endif


endmodule // OR5HSX4
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:44 and Version :1.1 //
 
//  START 
// CELL OR6HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR6HS_F_F_Z_F 0.1
`define OR6HS_F_R_Z_R 0.1
`define OR6HS_E_F_Z_F 0.1
`define OR6HS_E_R_Z_R 0.1
`define OR6HS_D_F_Z_F 0.1
`define OR6HS_D_R_Z_R 0.1
`define OR6HS_C_F_Z_F 0.1
`define OR6HS_C_R_Z_R 0.1
`define OR6HS_B_F_Z_F 0.1
`define OR6HS_B_R_Z_R 0.1
`define OR6HS_A_F_Z_F 0.1
`define OR6HS_A_R_Z_R 0.1

module OR6HS (Z, A, B, C, D, E, F);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;


   or  u0 (Z, A, B, C, D, E, F);


`ifdef functional
`else
   specify

      (F +=> Z) = (`OR6HS_F_R_Z_R,`OR6HS_F_F_Z_F);
      (E +=> Z) = (`OR6HS_E_R_Z_R,`OR6HS_E_F_Z_F);
      (D +=> Z) = (`OR6HS_D_R_Z_R,`OR6HS_D_F_Z_F);
      (C +=> Z) = (`OR6HS_C_R_Z_R,`OR6HS_C_F_Z_F);
      (B +=> Z) = (`OR6HS_B_R_Z_R,`OR6HS_B_F_Z_F);
      (A +=> Z) = (`OR6HS_A_R_Z_R,`OR6HS_A_F_Z_F);

   endspecify
`endif


endmodule // OR6HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:20:54 and Version :1.1 //
 
//  START 
// CELL OR7HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR7HS_G_F_Z_F 0.1
`define OR7HS_G_R_Z_R 0.1
`define OR7HS_F_F_Z_F 0.1
`define OR7HS_F_R_Z_R 0.1
`define OR7HS_E_F_Z_F 0.1
`define OR7HS_E_R_Z_R 0.1
`define OR7HS_D_F_Z_F 0.1
`define OR7HS_D_R_Z_R 0.1
`define OR7HS_C_F_Z_F 0.1
`define OR7HS_C_R_Z_R 0.1
`define OR7HS_B_F_Z_F 0.1
`define OR7HS_B_R_Z_R 0.1
`define OR7HS_A_F_Z_F 0.1
`define OR7HS_A_R_Z_R 0.1

module OR7HS (Z, A, B, C, D, E, F, G);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;
   input G;


   or  u0 (Z, A, B, C, D, E, F, G);


`ifdef functional
`else
   specify

      (G +=> Z) = (`OR7HS_G_R_Z_R,`OR7HS_G_F_Z_F);
      (F +=> Z) = (`OR7HS_F_R_Z_R,`OR7HS_F_F_Z_F);
      (E +=> Z) = (`OR7HS_E_R_Z_R,`OR7HS_E_F_Z_F);
      (D +=> Z) = (`OR7HS_D_R_Z_R,`OR7HS_D_F_Z_F);
      (C +=> Z) = (`OR7HS_C_R_Z_R,`OR7HS_C_F_Z_F);
      (B +=> Z) = (`OR7HS_B_R_Z_R,`OR7HS_B_F_Z_F);
      (A +=> Z) = (`OR7HS_A_R_Z_R,`OR7HS_A_F_Z_F);

   endspecify
`endif


endmodule // OR7HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:21:00 and Version :1.1 //
 
//  START 
// CELL OR8HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define OR8HS_H_F_Z_F 0.1
`define OR8HS_H_R_Z_R 0.1
`define OR8HS_G_F_Z_F 0.1
`define OR8HS_G_R_Z_R 0.1
`define OR8HS_F_F_Z_F 0.1
`define OR8HS_F_R_Z_R 0.1
`define OR8HS_E_F_Z_F 0.1
`define OR8HS_E_R_Z_R 0.1
`define OR8HS_D_F_Z_F 0.1
`define OR8HS_D_R_Z_R 0.1
`define OR8HS_C_F_Z_F 0.1
`define OR8HS_C_R_Z_R 0.1
`define OR8HS_B_F_Z_F 0.1
`define OR8HS_B_R_Z_R 0.1
`define OR8HS_A_F_Z_F 0.1
`define OR8HS_A_R_Z_R 0.1

module OR8HS (Z, A, B, C, D, E, F, G, H);

   output Z;
   input A;
   input B;
   input C;
   input D;
   input E;
   input F;
   input G;
   input H;


   or  u0 (Z, A, B, C, D, E, F, G, H);


`ifdef functional
`else
   specify

      (H +=> Z) = (`OR8HS_H_R_Z_R,`OR8HS_H_F_Z_F);
      (G +=> Z) = (`OR8HS_G_R_Z_R,`OR8HS_G_F_Z_F);
      (F +=> Z) = (`OR8HS_F_R_Z_R,`OR8HS_F_F_Z_F);
      (E +=> Z) = (`OR8HS_E_R_Z_R,`OR8HS_E_F_Z_F);
      (D +=> Z) = (`OR8HS_D_R_Z_R,`OR8HS_D_F_Z_F);
      (C +=> Z) = (`OR8HS_C_R_Z_R,`OR8HS_C_F_Z_F);
      (B +=> Z) = (`OR8HS_B_R_Z_R,`OR8HS_B_F_Z_F);
      (A +=> Z) = (`OR8HS_A_R_Z_R,`OR8HS_A_F_Z_F);

   endspecify
`endif


endmodule // OR8HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:21:06 and Version :1.1 //
 
//  END
// Created from CVS on Date :1998/07/08 13:43:50 and Version :1.3 //
 
//  START 
// CELL SCBTNBHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define SCBTNBHS_SD_F_CO_R 0.1
`define SCBTNBHS_CD_F_CO_F 0.1
`define SCBTNBHS_CD_R_CO_R 0.1
`define SCBTNBHS_CP_R_CO_F 0.1
`define SCBTNBHS_CP_R_CO_R 0.1
`define SCBTNBHS_CI_F_CO_F 0.1
`define SCBTNBHS_CI_R_CO_R 0.1
`define SCBTNBHS_SD_F_QN_F 0.1
`define SCBTNBHS_CD_F_QN_R 0.1
`define SCBTNBHS_CD_R_QN_F 0.1
`define SCBTNBHS_CP_R_QN_R 0.1
`define SCBTNBHS_CP_R_QN_F 0.1
`define SCBTNBHS_SD_F_Q_R 0.1
`define SCBTNBHS_CD_F_Q_F 0.1
`define SCBTNBHS_CD_R_Q_R 0.1
`define SCBTNBHS_CP_R_Q_F 0.1
`define SCBTNBHS_CP_R_Q_R 0.1
`define SCBTNBHS_CI_CP_HOLD_negedge_posedge 0.1
`define SCBTNBHS_CI_CP_SETUP_posedge_posedge 0.1
`define SCBTNBHS_CI_CP_HOLD_posedge_posedge 0.1
`define SCBTNBHS_CI_CP_SETUP_negedge_posedge 0.1
`define SCBTNBHS_CP_PWL 0.1
`define SCBTNBHS_CP_PWH 0.1
`define SCBTNBHS_SD_PWL 0.1
`define SCBTNBHS_CD_PWL 0.1
`define SCBTNBHS_SD_CP_REC_posedge_posedge 0.1
`define SCBTNBHS_CD_CP_REC_posedge_posedge 0.1
`define SCBTNBHS_SD_CP_REM_posedge_posedge 0.1
`define SCBTNBHS_CD_CP_REM_posedge_posedge 0.1
`define SCBTNBHS_CD_SD_REC_posedge_posedge 0.1
`define SCBTNBHS_CD_SD_REM_posedge_posedge 0.1

module SCBTNBHS (Q, QN, CO, CI, CP, CD, SD);

   output Q;
   output QN;
   output CO;
   input CI;
   input CP;
   input CD;
   input SD;


   reg Notifier;

   xor  u0 (XorCIIQ_, CI, IQ);

   U_FD_P_RN_SN_NOTI u1 (IQ, XorCIIQ_, CP, CD, SD, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);
   and  u4 (CO, CI, IQ);



`ifdef functional
`else
   and  (AndCDSD_, CD, SD);
   specify
`ifdef verifault

      (CI +=> CO) = (`SCBTNBHS_CI_R_CO_R,`SCBTNBHS_CI_F_CO_F);
      if(!IQ && CD && SD) (posedge CP => (Q +: CI)) = (`SCBTNBHS_CP_R_Q_R, `SCBTNBHS_CP_R_Q_F);
      if(IQ && CD && SD) (posedge CP => (Q -: CI)) = (`SCBTNBHS_CP_R_Q_R, `SCBTNBHS_CP_R_Q_F);
      if(!IQ && CD && SD) (posedge CP => (QN -: CI)) = (`SCBTNBHS_CP_R_QN_R, `SCBTNBHS_CP_R_QN_F);
      if(IQ && CD && SD) (posedge CP => (QN +: CI)) = (`SCBTNBHS_CP_R_QN_R, `SCBTNBHS_CP_R_QN_F);
      if(CI && CD && SD) (posedge CP => (CO +: IQ)) = (`SCBTNBHS_CP_R_CO_R, `SCBTNBHS_CP_R_CO_F);
      if(!SD) (posedge CD => (Q +: 1'b1)) = (`SCBTNBHS_CD_R_Q_R,`SCBTNBHS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`SCBTNBHS_CD_R_Q_R,`SCBTNBHS_CD_F_Q_F);
      if(CD) (negedge SD => (Q +: 1'b1)) = (`SCBTNBHS_SD_F_Q_R,`SCBTNBHS_SD_F_Q_R);
      if(!SD) (posedge CD => (QN +: 1'b0)) = (`SCBTNBHS_CD_F_QN_R,`SCBTNBHS_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`SCBTNBHS_CD_F_QN_R,`SCBTNBHS_CD_R_QN_F);
      if(CD) (negedge SD => (QN +: 1'b0)) = (`SCBTNBHS_SD_F_QN_F,`SCBTNBHS_SD_F_QN_F);
      if(CI && !SD) (posedge CD => (CO +: 1'b1)) = (`SCBTNBHS_CD_R_CO_R,`SCBTNBHS_CD_F_CO_F);
      (negedge CD => (CO +: 1'b0)) = (`SCBTNBHS_CD_R_CO_R,`SCBTNBHS_CD_F_CO_F);
      if(CI && CD) (negedge SD => (CO +: 1'b1)) = (`SCBTNBHS_SD_F_CO_R,`SCBTNBHS_SD_F_CO_R);

	$setuphold(posedge CP &&& AndCDSD_, posedge CI, `SCBTNBHS_CI_CP_SETUP_posedge_posedge, `SCBTNBHS_CI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& AndCDSD_, negedge CI, `SCBTNBHS_CI_CP_SETUP_negedge_posedge, `SCBTNBHS_CI_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `SCBTNBHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `SCBTNBHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `SCBTNBHS_SD_PWL, 0, Notifier);
      $width(negedge CD, `SCBTNBHS_CD_PWL, 0, Notifier);
	$recovery(posedge SD, posedge CP &&& CD, `SCBTNBHS_SD_CP_REC_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge CP &&& SD, `SCBTNBHS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP &&& CD, posedge SD, `SCBTNBHS_SD_CP_REM_posedge_posedge, Notifier);

	$hold(posedge CP &&& SD, posedge CD, `SCBTNBHS_CD_CP_REM_posedge_posedge, Notifier);

	$recovery(posedge CD, posedge SD, `SCBTNBHS_CD_SD_REC_posedge_posedge, Notifier);

	$hold(posedge SD, posedge CD, `SCBTNBHS_CD_SD_REM_posedge_posedge, Notifier);
`else

      (CI +=> CO) = (`SCBTNBHS_CI_R_CO_R,`SCBTNBHS_CI_F_CO_F);
      (posedge CP => (Q +: CI)) = (`SCBTNBHS_CP_R_Q_R, `SCBTNBHS_CP_R_Q_F);
      (posedge CP => (QN -: CI)) = (`SCBTNBHS_CP_R_QN_R, `SCBTNBHS_CP_R_QN_F);
      (posedge CP => (CO +: IQ)) = (`SCBTNBHS_CP_R_CO_R, `SCBTNBHS_CP_R_CO_F);
      (posedge CD => (Q +: 1'b1)) = (`SCBTNBHS_CD_R_Q_R,`SCBTNBHS_CD_F_Q_F);
      (negedge CD => (Q +: 1'b0)) = (`SCBTNBHS_CD_R_Q_R,`SCBTNBHS_CD_F_Q_F);
      (negedge SD => (Q +: 1'b1)) = (`SCBTNBHS_SD_F_Q_R,`SCBTNBHS_SD_F_Q_R);
      (posedge CD => (QN +: 1'b0)) = (`SCBTNBHS_CD_F_QN_R,`SCBTNBHS_CD_R_QN_F);
      (negedge CD => (QN +: 1'b1)) = (`SCBTNBHS_CD_F_QN_R,`SCBTNBHS_CD_R_QN_F);
      (negedge SD => (QN +: 1'b0)) = (`SCBTNBHS_SD_F_QN_F,`SCBTNBHS_SD_F_QN_F);
      (posedge CD => (CO +: 1'b1)) = (`SCBTNBHS_CD_R_CO_R,`SCBTNBHS_CD_F_CO_F);
      (negedge CD => (CO +: 1'b0)) = (`SCBTNBHS_CD_R_CO_R,`SCBTNBHS_CD_F_CO_F);
      (negedge SD => (CO +: 1'b1)) = (`SCBTNBHS_SD_F_CO_R,`SCBTNBHS_SD_F_CO_R);
 
        $setuphold(posedge CP &&& AndCDSD_, posedge CI, `SCBTNBHS_CI_CP_SETUP_posedge_posedge, `SCBTNBHS_CI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& AndCDSD_, negedge CI, `SCBTNBHS_CI_CP_SETUP_negedge_posedge, `SCBTNBHS_CI_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `SCBTNBHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& AndCDSD_, `SCBTNBHS_CP_PWH, 0, Notifier);
      $width(negedge SD, `SCBTNBHS_SD_PWL, 0, Notifier);
      $width(negedge CD, `SCBTNBHS_CD_PWL, 0, Notifier);
        $recovery(posedge SD, posedge CP &&& CD, `SCBTNBHS_SD_CP_REC_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge CP &&& SD, `SCBTNBHS_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& CD, posedge SD, `SCBTNBHS_SD_CP_REM_posedge_posedge, Notifier);
 
        $hold(posedge CP &&& SD, posedge CD, `SCBTNBHS_CD_CP_REM_posedge_posedge, Notifier);
 
        $recovery(posedge CD, posedge SD, `SCBTNBHS_CD_SD_REC_posedge_posedge, Notifier);
 
        $hold(posedge SD, posedge CD, `SCBTNBHS_CD_SD_REM_posedge_posedge, Notifier);
`endif

   endspecify
`endif


endmodule // SCBTNBHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/07 13:21:12 and Version :1.1 //
 
//  START 
// CELL SCCTNBHS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_unit
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define SCCTNBHS_CD_F_CO_F 0.1
`define SCCTNBHS_CP_R_CO_F 0.1
`define SCCTNBHS_CP_R_CO_R 0.1
`define SCCTNBHS_CI_F_CO_F 0.1
`define SCCTNBHS_CI_R_CO_R 0.1
`define SCCTNBHS_CD_F_QN_R 0.1
`define SCCTNBHS_CP_R_QN_R 0.1
`define SCCTNBHS_CP_R_QN_F 0.1
`define SCCTNBHS_CD_F_Q_F 0.1
`define SCCTNBHS_CP_R_Q_F 0.1
`define SCCTNBHS_CP_R_Q_R 0.1
`define SCCTNBHS_CI_CP_HOLD_negedge_posedge 0.1
`define SCCTNBHS_CI_CP_SETUP_posedge_posedge 0.1
`define SCCTNBHS_CI_CP_HOLD_posedge_posedge 0.1
`define SCCTNBHS_CI_CP_SETUP_negedge_posedge 0.1
`define SCCTNBHS_CP_PWL 0.1
`define SCCTNBHS_CP_PWH 0.1
`define SCCTNBHS_CD_PWL 0.1
`define SCCTNBHS_CD_CP_REC_posedge_posedge 0.1
`define SCCTNBHS_CD_CP_REM_posedge_posedge 0.1

module SCCTNBHS (Q, QN, CO, CI, CP, CD);

   output Q;
   output QN;
   output CO;
   input CI;
   input CP;
   input CD;


   reg Notifier;

   xor  u0 (XorCIIQ_, CI, IQ);

   U_FD_P_RN_NOTI u1 (IQ, XorCIIQ_, CP, CD, Notifier);

   buf  u2 (Q, IQ);
   not  u3 (QN, IQ);
   and  u4 (CO, CI, IQ);



`ifdef functional
`else
   specify
`ifdef verifault

      (CI +=> CO) = (`SCCTNBHS_CI_R_CO_R,`SCCTNBHS_CI_F_CO_F);
      if(!IQ && CD) (posedge CP => (Q +: CI)) = (`SCCTNBHS_CP_R_Q_R, `SCCTNBHS_CP_R_Q_F);
      if(IQ && CD) (posedge CP => (Q -: CI)) = (`SCCTNBHS_CP_R_Q_R, `SCCTNBHS_CP_R_Q_F);
      if(!IQ && CD) (posedge CP => (QN -: CI)) = (`SCCTNBHS_CP_R_QN_R, `SCCTNBHS_CP_R_QN_F);
      if(IQ && CD) (posedge CP => (QN +: CI)) = (`SCCTNBHS_CP_R_QN_R, `SCCTNBHS_CP_R_QN_F);
      if(CI && CD) (posedge CP => (CO +: IQ)) = (`SCCTNBHS_CP_R_CO_R, `SCCTNBHS_CP_R_CO_F);
      (negedge CD => (Q +: 1'b0)) = (`SCCTNBHS_CD_F_Q_F,`SCCTNBHS_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`SCCTNBHS_CD_F_QN_R,`SCCTNBHS_CD_F_QN_R);
      (negedge CD => (CO +: 1'b0)) = (`SCCTNBHS_CD_F_CO_F,`SCCTNBHS_CD_F_CO_F);

	$setuphold(posedge CP &&& CD, posedge CI, `SCCTNBHS_CI_CP_SETUP_posedge_posedge, `SCCTNBHS_CI_CP_HOLD_posedge_posedge, Notifier);
	$setuphold(posedge CP &&& CD, negedge CI, `SCCTNBHS_CI_CP_SETUP_negedge_posedge, `SCCTNBHS_CI_CP_HOLD_negedge_posedge, Notifier);

      $width(negedge CP, `SCCTNBHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `SCCTNBHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `SCCTNBHS_CD_PWL, 0, Notifier);
	$recovery(posedge CD, posedge CP, `SCCTNBHS_CD_CP_REC_posedge_posedge, Notifier);

	$hold(posedge CP, posedge CD, `SCCTNBHS_CD_CP_REM_posedge_posedge, Notifier);
`else

      (CI +=> CO) = (`SCCTNBHS_CI_R_CO_R,`SCCTNBHS_CI_F_CO_F);
      (posedge CP => (Q +: CI)) = (`SCCTNBHS_CP_R_Q_R, `SCCTNBHS_CP_R_Q_F);
      (posedge CP => (QN -: CI)) = (`SCCTNBHS_CP_R_QN_R, `SCCTNBHS_CP_R_QN_F);
      (posedge CP => (CO +: IQ)) = (`SCCTNBHS_CP_R_CO_R, `SCCTNBHS_CP_R_CO_F);
      (negedge CD => (Q +: 1'b0)) = (`SCCTNBHS_CD_F_Q_F,`SCCTNBHS_CD_F_Q_F);
      (negedge CD => (QN +: 1'b1)) = (`SCCTNBHS_CD_F_QN_R,`SCCTNBHS_CD_F_QN_R);
      (negedge CD => (CO +: 1'b0)) = (`SCCTNBHS_CD_F_CO_F,`SCCTNBHS_CD_F_CO_F);
 
        $setuphold(posedge CP &&& CD, posedge CI, `SCCTNBHS_CI_CP_SETUP_posedge_posedge, `SCCTNBHS_CI_CP_HOLD_posedge_posedge, Notifier);
        $setuphold(posedge CP &&& CD, negedge CI, `SCCTNBHS_CI_CP_SETUP_negedge_posedge, `SCCTNBHS_CI_CP_HOLD_negedge_posedge, Notifier);
 
      $width(negedge CP, `SCCTNBHS_CP_PWL, 0, Notifier);
      $width(posedge CP &&& CD, `SCCTNBHS_CP_PWH, 0, Notifier);
      $width(negedge CD, `SCCTNBHS_CD_PWL, 0, Notifier);
        $recovery(posedge CD, posedge CP, `SCCTNBHS_CD_CP_REC_posedge_posedge, Notifier);
 
        $hold(posedge CP, posedge CD, `SCCTNBHS_CD_CP_REM_posedge_posedge, Notifier);
`endif

   endspecify
`endif


endmodule // SCCTNBHS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END
// Created from CVS on Date :1998/07/08 13:43:50 and Version :1.3 //
 
//  START 
// CELL SU1HS

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define SU1HS_CI_F_CO_F 0.1
`define SU1HS_CI_R_CO_R 0.1
`define SU1HS_B_F_CO_R 0.1
`define SU1HS_B_R_CO_F 0.1
`define SU1HS_A_F_CO_F 0.1
`define SU1HS_A_R_CO_R 0.1
`define SU1HS_CI_F_Z_R 0.1
`define SU1HS_CI_R_Z_F 0.1
`define SU1HS_CI_F_Z_F 0.1
`define SU1HS_CI_R_Z_R 0.1
`define SU1HS_B_F_Z_R 0.1
`define SU1HS_B_R_Z_F 0.1
`define SU1HS_B_F_Z_F 0.1
`define SU1HS_B_R_Z_R 0.1
`define SU1HS_A_F_Z_R 0.1
`define SU1HS_A_R_Z_F 0.1
`define SU1HS_A_F_Z_F 0.1
`define SU1HS_A_R_Z_R 0.1

module SU1HS (Z, CO, A, B, CI);

   output Z;
   output CO;
   input A;
   input B;
   input CI;


   xnor  u0 (Z, A, B, CI);
   not  u1 (BX, B);
   or  u2 (OrABX_, A, BX);
   and  u3 (AndOrABX_CI_, OrABX_, CI);
   and  u4 (AndABX_, A, BX);
   or  u5 (CO, AndOrABX_CI_, AndABX_);


`ifdef functional
`else
   specify

      (CI +=> CO) = (`SU1HS_CI_R_CO_R,`SU1HS_CI_F_CO_F);
      (B -=> CO) = (`SU1HS_B_F_CO_R,`SU1HS_B_R_CO_F);
      (A +=> CO) = (`SU1HS_A_R_CO_R,`SU1HS_A_F_CO_F);
      if (A && B || !A && !B) (CI -=> Z) = (`SU1HS_CI_F_Z_R,`SU1HS_CI_R_Z_F);
      if (!A && B || A && !B) (CI +=> Z) = (`SU1HS_CI_R_Z_R,`SU1HS_CI_F_Z_F);
      if (A && CI || !A && !CI) (B -=> Z) = (`SU1HS_B_F_Z_R,`SU1HS_B_R_Z_F);
      if (!A && CI || A && !CI) (B +=> Z) = (`SU1HS_B_R_Z_R,`SU1HS_B_F_Z_F);
      if (B && CI || !B && !CI) (A -=> Z) = (`SU1HS_A_F_Z_R,`SU1HS_A_R_Z_F);
      if (!B && CI || B && !CI) (A +=> Z) = (`SU1HS_A_R_Z_R,`SU1HS_A_F_Z_F);

   endspecify
`endif


endmodule // SU1HS
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END

//  START
// CELL SU1HSP

`celldefine
`ifdef verifault
`suppress_faults
`enable_portfaults
`endif
`ifdef functional
   `timescale 1ns / 1ns
   `delay_mode_zero
`else
   `timescale 1ns / 10ps
   `delay_mode_path
`endif
 

`define SU1HSP_CI_F_CO_F 0.1
`define SU1HSP_CI_R_CO_R 0.1
`define SU1HSP_B_F_CO_R 0.1
`define SU1HSP_B_R_CO_F 0.1
`define SU1HSP_A_F_CO_F 0.1
`define SU1HSP_A_R_CO_R 0.1
`define SU1HSP_CI_F_Z_R 0.1
`define SU1HSP_CI_R_Z_F 0.1
`define SU1HSP_CI_F_Z_F 0.1
`define SU1HSP_CI_R_Z_R 0.1
`define SU1HSP_B_F_Z_R 0.1
`define SU1HSP_B_R_Z_F 0.1
`define SU1HSP_B_F_Z_F 0.1
`define SU1HSP_B_R_Z_R 0.1
`define SU1HSP_A_F_Z_R 0.1
`define SU1HSP_A_R_Z_F 0.1
`define SU1HSP_A_F_Z_F 0.1
`define SU1HSP_A_R_Z_R 0.1

module SU1HSP (Z, CO, A, B, CI);

   output Z;
   output CO;
   input A;
   input B;
   input CI;


   xnor  u0 (Z, A, B, CI);
   not  u1 (BX, B);
   or  u2 (OrABX_, A, BX);
   and  u3 (AndOrABX_CI_, OrABX_, CI);
   and  u4 (AndABX_, A, BX);
   or  u5 (CO, AndOrABX_CI_, AndABX_);


`ifdef functional
`else
   specify

      (CI +=> CO) = (`SU1HSP_CI_R_CO_R,`SU1HSP_CI_F_CO_F);
      (B -=> CO) = (`SU1HSP_B_F_CO_R,`SU1HSP_B_R_CO_F);
      (A +=> CO) = (`SU1HSP_A_R_CO_R,`SU1HSP_A_F_CO_F);
      if (A && B || !A && !B) (CI -=> Z) = (`SU1HSP_CI_F_Z_R,`SU1HSP_CI_R_Z_F);
      if (!A && B || A && !B) (CI +=> Z) = (`SU1HSP_CI_R_Z_R,`SU1HSP_CI_F_Z_F);
      if (A && CI || !A && !CI) (B -=> Z) = (`SU1HSP_B_F_Z_R,`SU1HSP_B_R_Z_F);
      if (!A && CI || A && !CI) (B +=> Z) = (`SU1HSP_B_R_Z_R,`SU1HSP_B_F_Z_F);
      if (B && CI || !B && !CI) (A -=> Z) = (`SU1HSP_A_F_Z_R,`SU1HSP_A_R_Z_F);
      if (!B && CI || B && !CI) (A +=> Z) = (`SU1HSP_A_R_Z_R,`SU1HSP_A_F_Z_F);

   endspecify
`endif


endmodule // SU1HSP
`ifdef verifault
`disable_portfaults
`nosuppress_faults
`endif
`endcelldefine


//  END

//  START


primitive U_FD_P_NOTI (Q, D, CP, NOTI_REG);

   output Q;
   input  D,		// data
          CP,		// clock
          NOTI_REG;
   reg    Q;

   table

      // D     CP    NOTI_REG    : Qtn : Qtn+1

         0     (01)  ?           :  ?  :  0  ;		// Normal clocking
         1     (01)  ?           :  ?  :  1  ;

         *     b     ?           :  ?  :  -  ;		// Ignore edges on data

         ?     (?0)  ?           :  ?  :  -  ;		// Ignore falling edges on clock

         0     (1x)  ?           :  0  :  0  ;		// Cases reducing pessimism
         1     (1x)  ?           :  1  :  1  ;
         0     (0x)  ?           :  0  :  0  ;
         0     (x1)  ?           :  0  :  0  ;
         1     (0x)  ?           :  1  :  1  ;
         1     (x1)  ?           :  1  :  1  ;

         ?     ?     *           :  ?  :  x  ;		// X for timing violations

   endtable

endprimitive


primitive U_FD_P_RN_NOTI (Q, D, CP, RN, NOTI_REG);

   output Q;
   input  D,		// data
          CP,		// clock
          RN,		// clear active low
          NOTI_REG;
   reg    Q;

   table
 
      // D     CP    RN    NOTI_REG    : Qtn : Qtn+1

         ?     ?     0     ?           :  ?  :  0  ;	// Asynchronous clear

         1     (01)  1     ?           :  ?  :  1  ;	// Normal clocking
         0     (01)  1     ?           :  ?  :  0  ;

         *     b     ?     ?           :  ?  :  -  ;	// Ignore edges on data

         ?     (?0)  ?     ?           :  ?  :  -  ;	// Ignore falling edges on clock

         0     (1x)  ?     ?           :  0  :  0  ;
         1     (1x)  1     ?           :  1  :  1  ;

         ?     b     (?1)  ?           :  ?  :  -  ;	// Ignore rising edges on clear
         0     x     (?1)  ?           :  0  :  0  ;	// Ignore rising edges on clear

         0     (0x)  ?     ?           :  0  :  0  ;	// Cases reducing pessimism
         0     (x1)  ?     ?           :  0  :  0  ;
         1     (0x)  1     ?           :  1  :  1  ;
         1     (x1)  1     ?           :  1  :  1  ;

         0     (01)  x     ?           :  ?  :  0  ;
         ?     b     (?x)  ?           :  0  :  0  ;
         0     x     (?x)  ?           :  0  :  0  ;

         ?     ?     ?     *           :  ?  :  x  ;	// X for timing violations

   endtable

endprimitive


primitive U_FD_P_RN_SN_NOTI (Q, D, CP, RN, SN, NOTI_REG);

   output Q;
   input  D,		// data
          CP,		// clock
          RN,		// clear active low
          SN,		// preset active low
          NOTI_REG;
   reg    Q;

   table

      // D     CP    RN    SN    NOTI_REG    : Qtn : Qtn+1

         ?     ?     0     ?     ?           :  ?  :  0  ;	// Asynchronous clear
         ?     ?     1     0     ?           :  ?  :  1  ;	// Asynchronous preset

         0     (01)  1     1     ?           :  ?  :  0  ;	// Normal clocking
         1     (01)  1     1     ?           :  ?  :  1  ;

         *     b     ?     ?     ?           :  ?  :  -  ;	// Ignore edges on data

         ?     (?0)  ?     ?     ?           :  ?  :  -  ;	// Ignore falling edges on clock
         1     (1x)  1     ?     ?           :  1  :  1  ;
         0     (1x)  ?     1     ?           :  0  :  0  ;

         ?     b     (?1)  1     ?           :  ?  :  -  ;	// Ignore rising edges on clear
         0     x     (?1)  1     ?           :  0  :  0  ;	// Ignore rising edges on clear
         ?     b     1     (?1)  ?           :  ?  :  -  ;	// Ignore rising edges on preset
         1     x     1     (?1)  ?           :  1  :  1  ;	// Ignore rising edges on preset

         0     (0x)  ?     1     ?           :  0  :  0  ;	// Cases reducing pessimism
         0     (x1)  ?     1     ?           :  0  :  0  ;
         1     (0x)  1     ?     ?           :  1  :  1  ;
         1     (x1)  1     ?     ?           :  1  :  1  ;

         0     (01)  x     1     ?           :  ?  :  0  ;
         ?     b     (?x)  1     ?           :  0  :  0  ;
         0     x     (?x)  1     ?           :  0  :  0  ;	// Line added

         1     (01)  1     x     ?           :  ?  :  1  ;
         ?     b     1     (?x)  ?           :  1  :  1  ;
         1     x     1     (?x)  ?           :  1  :  1  ;	// Line added

         ?     ?     ?     ?     *           :  ?  :  x  ;	// X for timing violations

   endtable

endprimitive


primitive U_FD_P_SN_NOTI (Q, D, CP, SN, NOTI_REG);

   output Q;
   input  D,		// data
          CP,		// clock
          SN,		// preset active low
          NOTI_REG;
   reg    Q;

   table
 
      // D     CP    SN    NOTI_REG    : Qtn : Qtn+1

         ?     ?     0     ?           :  ?  :  1  ;	// Asynchronous preset

         1     (01)  1     ?           :  ?  :  1  ;	// Normal clocking
         0     (01)  1     ?           :  ?  :  0  ;

         *     b     ?     ?           :  ?  :  -  ;	// Ignore edges on data

         ?     (?0)  ?     ?           :  ?  :  -  ;	// Ignore falling edges on clock

         0     (1x)  1     ?           :  0  :  0  ;
         1     (1x)  ?     ?           :  1  :  1  ;

         ?     b     (?1)  ?           :  ?  :  -  ;	// Ignore rising edges on set
         1     x     (?1)  ?           :  1  :  1  ;	// Ignore rising edges on set

         0     (0x)  1     ?           :  0  :  0  ;	// Cases reducing pessimism
         0     (x1)  1     ?           :  0  :  0  ;
         1     (0x)  ?     ?           :  1  :  1  ;
         1     (x1)  ?     ?           :  1  :  1  ;

         1     (01)  x     ?           :  ?  :  1  ;
         ?     b     (?x)  ?           :  1  :  1  ;
         1     x     (?x)  ?           :  1  :  1  ;

         ?     ?     ?     *           :  ?  :  x  ;	// X for timing violations

   endtable

endprimitive


primitive U_LD_N_NOTI (Q, D, GN, NOTI_REG);
 
   output Q;
   input  D,            // data
          GN,           // clock active low
          NOTI_REG;
   reg    Q;
 
   table
 
      // D     GN    NOTI_REG    : Qtn : Qtn+1
 
         (?0)  0     ?           :  ?  :  0  ;          // Transparency
         (?1)  0     ?           :  ?  :  1  ;
 
         0     (?0)  ?           :  ?  :  0  ;
         1     (?0)  ?           :  ?  :  1  ;
 
         *     1     ?           :  ?  :  -  ;          // Latching
 
         ?     (?1)  ?           :  ?  :  -  ;          // Ignore rising edges on clock
         ?     (0x)  ?           :  ?  :  -  ;
 
         0     (1x)  ?           :  0  :  0  ;          // Cases reducing pessimism
         1     (1x)  ?           :  1  :  1  ;
         (?0)  x     ?           :  0  :  0  ;
         (?1)  x     ?           :  1  :  1  ;
 
         ?     ?     *           :  ?  :  x  ;          // X for timing violations
 
   endtable
 

endprimitive


primitive U_LD_N_RN_NOTI (Q, D, GN, RN, NOTI_REG);
 
   output Q;
   input  D,            // data
          GN,           // clock active low
          RN,           // clear active low
          NOTI_REG;
   reg    Q;
 
   table
 
      // D     GN    RN    NOTI_REG : Qtn : Qtn+1
 
         ?     ?     0     ?        :  ?  :  0  ;       // Asynchronous clear
 
         (?0)  0     1     ?        :  ?  :  0  ;       // Transparency
         (?1)  0     1     ?        :  ?  :  1  ;
 
         0     (?0)  1     ?        :  ?  :  0  ;
         1     (?0)  1     ?        :  ?  :  1  ;
 
         *     1     1     ?        :  ?  :  -  ;       // Latching
         *     1     x     ?        :  ?  :  -  ;
 
         ?     (?1)  ?     ?        :  ?  :  -  ;       // Ignore rising edges on clock
         ?     (0x)  ?     ?        :  ?  :  -  ;
 
         ?     1     (?1)  ?        :  ?  :  -  ;       // Rising edge on clear
         0     0     (?1)  ?        :  ?  :  0  ;
         1     0     (?1)  ?        :  ?  :  1  ;
         0     X     (?1)  ?        :  0  :  0  ;
 
         0     (1x)  1     ?        :  0  :  0  ;       // Cases reducing pessimism
         1     (1x)  1     ?        :  1  :  1  ;
         0     (1x)  X     ?        :  0  :  0  ;
 
         (?0)  x     1     ?        :  0  :  0  ;
         (?1)  x     1     ?        :  1  :  1  ;
 
         (?0)  0     x     ?        :  ?  :  0  ;
         0     (?0)  x     ?        :  ?  :  0  ;
 
         0     ?     (?x)  ?        :  0  :  0  ;
         1     1     (?x)  ?        :  0  :  0  ;
         X     1     (?x)  ?        :  0  :  0  ;
         ?     ?     ?     *        :  ?  :  x  ;       // X for timing violations

   endtable
 
endprimitive


primitive U_LD_N_RN_SN_NOTI (Q, D, GN, RN, SN, NOTI_REG);
 
   output Q;
   input  D,            // data
          GN,           // clock
          RN,           // clear active low
          SN,           // preset active low
          NOTI_REG;
   reg    Q;
 
   table
 
      // D     GN    RN    SN    NOTI_REG : Qtn : Qtn+1
 
         ?     ?     0     1     ?        :  ?  :  0  ; // Asynchronous clear
         ?     ?     ?     0     ?        :  ?  :  1  ; // Asynchronous preset
 
         (?0)  0     1     1     ?        :  ?  :  0  ; // Transparency
         (?1)  0     1     1     ?        :  ?  :  1  ;
 
         0     (?0)  1     1     ?        :  ?  :  0  ;
         1     (?0)  1     1     ?        :  ?  :  1  ;
 
         *     1     1     1     ?        :  ?  :  -  ; // Latching
         *     1     x     1     ?        :  ?  :  -  ;
         *     1     1     x     ?        :  ?  :  -  ;
 
         ?     (?1)  ?     ?     ?        :  ?  :  -  ; // Ignore rising edges on clock
         ?     (0x)  ?     ?     ?        :  ?  :  -  ;
 
         ?     1     (?1)  1     ?        :  ?  :  -  ; // Rising edge on clear
         0     0     (?1)  1     ?        :  ?  :  0  ;
         1     0     (?1)  1     ?        :  ?  :  1  ;
         1     0     (?1)  X     ?        :  ?  :  1  ;
         0     X     (?1)  1     ?        :  0  :  0  ;
 
         ?     1     1     (?1)  ?        :  ?  :  -  ; // Rising edge on preset
         0     0     1     (?1)  ?        :  ?  :  0  ;
         0     0     X     (?1)  ?        :  ?  :  0  ;
         1     0     1     (?1)  ?        :  ?  :  1  ;
         1     X     1     (?1)  ?        :  1  :  1  ;
 
         0     (1x)  1     1     ?        :  0  :  0  ; // Cases reducing pessimism
         0     (1x)  X     1     ?        :  0  :  0  ; // Cases reducing pessimism
         1     (1x)  1     1     ?        :  1  :  1  ;
         1     (1x)  1     X     ?        :  1  :  1  ;
         (?0)  x     1     1     ?        :  0  :  0  ;
         (?1)  x     1     1     ?        :  1  :  1  ;
 
         (?0)  0     x     1     ?        :  ?  :  0  ;
         0     (?0)  x     1     ?        :  ?  :  0  ;
 
         (?1)  0     1     x     ?        :  ?  :  1  ;
         1     (?0)  1     x     ?        :  ?  :  1  ;
 
//       ?     ?     (?x)  1     ?        :  0  :  0  ;
         0     ?     (?x)  1     ?        :  0  :  0  ;
         1     1     (?x)  1     ?        :  0  :  0  ;
         X     1     (?x)  1     ?        :  0  :  0  ;
 
//       ?     ?     1     (?x)  ?        :  1  :  1  ;
         1     ?     1     (?x)  ?        :  1  :  1  ;
         0     1     1     (?x)  ?        :  1  :  1  ;
         X     1     1     (?x)  ?        :  1  :  1  ;
 
         ?     ?     ?     ?     *        :  ?  :  x  ; // X for timing violations
 
   endtable
 
endprimitive


primitive U_LD_N_SN_NOTI (Q, D, GN, SN, NOTI_REG);
 
   output Q;
   input  D,            // data
          GN,           // clock
          SN,           // preset active low
          NOTI_REG;
   reg    Q;
 
   table
 
      // D     GN    SN    NOTI_REG : Qtn : Qtn+1
 
         ?     ?     0     ?        :  ?  :  1  ;       // Asynchronous preset
 
         (?0)  0     1     ?        :  ?  :  0  ;       // Transparency
         (?1)  0     1     ?        :  ?  :  1  ;
 
         0     (?0)  1     ?        :  ?  :  0  ;
         1     (?0)  1     ?        :  ?  :  1  ;
 
         *     1     1     ?        :  ?  :  -  ;       // Latching
         *     1     x     ?        :  ?  :  -  ;
 
         ?     (?1)  ?     ?        :  ?  :  -  ;       // Ignore rising edges on clock
         ?     (0x)  ?     ?        :  ?  :  -  ;
 
         ?     1     (?1)  ?        :  ?  :  -  ;       // Rising edge on preset
         0     0     (?1)  ?        :  ?  :  0  ;
         1     0     (?1)  ?        :  ?  :  1  ;
         1     X     (?1)  ?        :  1  :  1  ;
 
         0     (1x)  1     ?        :  0  :  0  ;       // Cases reducing pessimism
         1     (1x)  1     ?        :  1  :  1  ;
         1     (1x)  X     ?        :  1  :  1  ;
 
         (?0)  x     1     ?        :  0  :  0  ;
         (?1)  x     1     ?        :  1  :  1  ;
 
         (?1)  0     x     ?        :  ?  :  1  ;
         1     (?0)  x     ?        :  ?  :  1  ;
 
         1     ?     (?x)  ?        :  1  :  1  ;
         0     1     (?x)  ?        :  1  :  1  ;
         X     1     (?x)  ?        :  1  :  1  ;
         ?     ?     ?     *        :  ?  :  x  ;       // X for timing violations

   endtable
 
endprimitive


primitive U_LD_P_NOTI (Q, D, G, NOTI_REG);
 
   output Q;
   input  D,            // data
          G,            // clock
          NOTI_REG;
   reg    Q;
 
   table
 
      // D     G     NOTI_REG    : Qtn : Qtn+1
 
         (?0)  1     ?           :  ?  :  0  ;          // Transparency
         (?1)  1     ?           :  ?  :  1  ;
 
         0     (?1)  ?           :  ?  :  0  ;
         1     (?1)  ?           :  ?  :  1  ;
 
         *     0     ?           :  ?  :  -  ;          // Latching
 
         ?     (?0)  ?           :  ?  :  -  ;          // Ignore falling edges on clock
         ?     (1x)  ?           :  ?  :  -  ;
 
         0     (0x)  ?           :  0  :  0  ;          // Cases reducing pessimism
         1     (0x)  ?           :  1  :  1  ;
         (?0)  x     ?           :  0  :  0  ;
         (?1)  x     ?           :  1  :  1  ;
 
         ?     ?     *           :  ?  :  x  ;          // X for timing violations
 
   endtable
 

endprimitive


primitive U_LD_P_RN_NOTI (Q, D, G, RN, NOTI_REG);
 
   output Q;
   input  D,            // data
          G,            // clock
          RN,           // clear active low
          NOTI_REG;
   reg    Q;
 
   table
 
      // D     G     RN    NOTI_REG : Qtn : Qtn+1
 
         ?     ?     0     ?        :  ?  :  0  ;       // Asynchronous clear
 
         (?0)  1     1     ?        :  ?  :  0  ;       // Transparency
         (?1)  1     1     ?        :  ?  :  1  ;
 
         0     (?1)  1     ?        :  ?  :  0  ;
         1     (?1)  1     ?        :  ?  :  1  ;
 
         *     0     1     ?        :  ?  :  -  ;       // Latching
         *     0     x     ?        :  ?  :  -  ;
 
         ?     (?0)  ?     ?        :  ?  :  -  ;       // Ignore falling edges on clock
         ?     (1x)  ?     ?        :  ?  :  -  ;
 
         ?     0     (?1)  ?        :  ?  :  -  ;       // Rising edge on clear
         0     1     (?1)  ?        :  ?  :  0  ;
         1     1     (?1)  ?        :  ?  :  1  ;
         0     X     (?1)  ?        :  0  :  0  ;
 
         0     (0x)  1     ?        :  0  :  0  ;       // Cases reducing pessimism
         1     (0x)  1     ?        :  1  :  1  ;
         0     (0x)  X     ?        :  0  :  0  ;
 
         (?0)  x     1     ?        :  0  :  0  ;
         (?1)  x     1     ?        :  1  :  1  ;
 
         (?0)  1     x     ?        :  ?  :  0  ;
         0     (?1)  x     ?        :  ?  :  0  ;
 
         0     ?     (?x)  ?        :  0  :  0  ;
         1     0     (?x)  ?        :  0  :  0  ;
         X     0     (?x)  ?        :  0  :  0  ;
         ?     ?     ?     *        :  ?  :  x  ;       // X for timing violations

   endtable
 
endprimitive


primitive U_LD_P_SN_NOTI (Q, D, G, SN, NOTI_REG);
 
   output Q;
   input  D,            // data
          G,            // clock
          SN,           // preset active low
          NOTI_REG;
   reg    Q;
 
   table
 
      // D     G     SN    NOTI_REG : Qtn : Qtn+1
 
         ?     ?     0     ?        :  ?  :  1  ;       // Asynchronous preset
 
         (?0)  1     1     ?        :  ?  :  0  ;       // Transparency
         (?1)  1     1     ?        :  ?  :  1  ;
 
         0     (?1)  1     ?        :  ?  :  0  ;
         1     (?1)  1     ?        :  ?  :  1  ;
 
         *     0     1     ?        :  ?  :  -  ;       // Latching
         *     0     x     ?        :  ?  :  -  ;
 
         ?     (?0)  ?     ?        :  ?  :  -  ;       // Ignore falling edges on clock
         ?     (1x)  ?     ?        :  ?  :  -  ;
 
         ?     0     (?1)  ?        :  ?  :  -  ;       // Rising edge on preset
         0     1     (?1)  ?        :  ?  :  0  ;
         1     1     (?1)  ?        :  ?  :  1  ;
         1     X     (?1)  ?        :  1  :  1  ;
 
         0     (0x)  1     ?        :  0  :  0  ;       // Cases reducing pessimism
         1     (0x)  1     ?        :  1  :  1  ;
         1     (0x)  X     ?        :  1  :  1  ;
 
         (?0)  x     1     ?        :  0  :  0  ;
         (?1)  x     1     ?        :  1  :  1  ;
 
         (?1)  1     x     ?        :  ?  :  1  ;
         1     (?1)  x     ?        :  ?  :  1  ;
 
         1     ?     (?x)  ?        :  1  :  1  ;
         0     0     (?x)  ?        :  1  :  1  ;
         X     0     (?x)  ?        :  1  :  1  ;
         ?     ?     ?     *        :  ?  :  x  ;       // X for timing violations
 
   endtable
 
endprimitive


primitive U_MAJ (CO, A, B, CI);

   output CO;
   input A, B, CI;

   table

      // A  B  CI :  CO

         0  0  ?  :  0  ;
         0  ?  0  :  0  ;
         ?  0  0  :  0  ;
         1  1  ?  :  1  ;
         1  ?  1  :  1  ;
         ?  1  1  :  1  ;

   endtable

endprimitive


primitive U_MUX2 (Z, A, B, S);

   output Z;
   input  A, B, S;

   table

      // A  B  S  :  Z

         0  ?  0  :  0  ;
         1  ?  0  :  1  ;

         ?  0  1  :  0  ;
         ?  1  1  :  1  ;

      // Cases reducing pessimism

         0  0  x  :  0  ;
         1  1  x  :  1  ;

   endtable


endprimitive


primitive U_MUX4 (Y, D0, D1, D2, D3, S0, S1);

   output Y;
   input  D0, D1, D2, D3, S0, S1;

   table

      // D0 D1 D2 D3 S0 S1 :  Y

         0  ?  ?  ?  0  0  :  0  ;
         1  ?  ?  ?  0  0  :  1  ;

         ?  0  ?  ?  1  0  :  0  ;
         ?  1  ?  ?  1  0  :  1  ;

         ?  ?  0  ?  0  1  :  0  ;
         ?  ?  1  ?  0  1  :  1  ;

         ?  ?  ?  0  1  1  :  0  ;
         ?  ?  ?  1  1  1  :  1  ;

      // Cases reducing pessimism

         0  0  ?  ?  x  0  :  0  ;
         1  1  ?  ?  x  0  :  1  ;

         ?  ?  0  0  x  1  :  0  ;
         ?  ?  1  1  x  1  :  1  ;

         0  ?  0  ?  0  x  :  0  ;
         1  ?  1  ?  0  x  :  1  ;

         ?  0  ?  0  1  x  :  0  ;
         ?  1  ?  1  1  x  :  1  ;

         0  0  0  0  x  x  :  0  ;
         1  1  1  1  x  x  :  1  ;

   endtable

endprimitive


primitive U_RS_RN_SN_NOTI (Q, RN, SN, NOTI_REG);
 
   output Q;
   input  RN,            // reset
          SN,            // set
          NOTI_REG;
   reg    Q;
 
   table
 
      // RN     SN    NOTI_REG : Qtn : Qtn+1
         (?0)   ?        ?     :  ?  :  0  ;
         0      *        ?     :  ?  :  0  ;
         (?1)   0        ?     :  ?  :  1  ;
         1      (?0)     ?     :  ?  :  1  ;
 
         (?1)   1        ?     :  ?  :  -  ;
         1      (?1)     ?     :  ?  :  -  ;
 
         1      *        ?     :  1  :  1  ;
 
         *      1        ?     :  0  :  0  ;
 
         ?      ?        *     :  ?  :  x  ;       // X for timing violations
 
   endtable
 
 
endprimitive
