// SCHEMATIC SPICE SIM w/o EXTRACTION

module ring_gen100 (clk_out, rst_n);

	input  rst_n;
	output clk_out;

	wire rst_n;
	wire clok_out;

	wire w01i, w01o;
	wire w02i, w02o;
	wire w03i, w03o;
	wire w04i, w04o;
	wire w05i, w05o;
	wire w06i, w06o;
	wire w07i, w07o;
	wire w08i, w08o;
	wire w09i, w09o;
	wire w10i, w10o;
	wire w11i, w11o;
	wire w12i, w12o;
	wire w13i, w13o;
	wire w14i, w14o;
	wire w15i, w15o;
	wire w16i, w16o;
	wire w17i, w17o;
	wire w18i, w18o;
	wire w19i, w19o;
	wire w20i, w20o;
	wire w21i, w21o;
	wire w22i, w22o;
	wire w23i, w23o;
	wire w24i, w24o;
	wire w25i, w25o;
	wire w26i, w26o;
	wire w27i, w27o;
	wire w28i, w28o;
	wire w29i, w29o;
	wire w30i, w30o;
	wire w31i, w31o;
	wire w32i, w32o;
	wire w33i, w33o;
	wire w34i, w34o;
	wire w35i, w35o;
	wire w36i, w36o;
	wire w37i, w37o;
	wire w38i, w38o;
	wire w39i, w39o;
	wire w40i, w40o;
	wire w41i, w41o;
	wire w42i, w42o;
	wire w43i, w43o;
	wire w44i, w44o;
	wire w45i, w45o;
	wire w46i, w46o;
	wire w47i, w47o;
	wire w48i, w48o;
	wire w49i, w49o;
	wire w50i, w50o;
	wire w51i, w51o;
	wire w52i, w52o;
	wire w53i, w53o;

	wire wi, wo, diff_lb;

	IVHSP inv001 (.A(wi), .Z(w01o));
	IVHSP inv002 (.A(w01o), .Z(w02i));
	IVHSP inv003 (.A(w02i), .Z(w02o));
	IVHSP inv004 (.A(w02o), .Z(w03i));
	IVHSP inv005 (.A(w03i), .Z(w03o));
	IVHSP inv006 (.A(w03o), .Z(w04i));
	IVHSP inv007 (.A(w04i), .Z(w04o));
	IVHSP inv008 (.A(w04o), .Z(w05i));
	IVHSP inv009 (.A(w05i), .Z(w05o));
	IVHSP inv010 (.A(w05o), .Z(w06i));
	IVHSP inv011 (.A(w06i), .Z(w06o));
	IVHSP inv012 (.A(w06o), .Z(w07i));
	IVHSP inv013 (.A(w07i), .Z(w07o));
	IVHSP inv014 (.A(w07o), .Z(w08i));
	IVHSP inv015 (.A(w08i), .Z(w08o));
	IVHSP inv016 (.A(w08o), .Z(w09i));
	IVHSP inv017 (.A(w09i), .Z(w09o));
	IVHSP inv018 (.A(w09o), .Z(w10i));
	IVHSP inv019 (.A(w10i), .Z(w10o));
	IVHSP inv020 (.A(w10o), .Z(w11i));
	IVHSP inv021 (.A(w11i), .Z(w11o));
	IVHSP inv022 (.A(w11o), .Z(w12i));
	IVHSP inv023 (.A(w12i), .Z(w12o));
	IVHSP inv024 (.A(w12o), .Z(w13i));
	IVHSP inv025 (.A(w13i), .Z(w13o));
	IVHSP inv026 (.A(w13o), .Z(w14i));
	IVHSP inv027 (.A(w14i), .Z(w14o));
	IVHSP inv028 (.A(w14o), .Z(w15i));
	IVHSP inv029 (.A(w15i), .Z(w15o));
	IVHSP inv030 (.A(w15o), .Z(w16i));
	IVHSP inv031 (.A(w16i), .Z(w16o));
	IVHSP inv032 (.A(w16o), .Z(w17i));
	IVHSP inv033 (.A(w17i), .Z(w17o));
	IVHSP inv034 (.A(w17o), .Z(w18i));
	IVHSP inv035 (.A(w18i), .Z(w18o));
	IVHSP inv036 (.A(w18o), .Z(w19i));
	IVHSP inv037 (.A(w19i), .Z(w19o));
	IVHSP inv038 (.A(w19o), .Z(w20i));
	IVHSP inv039 (.A(w20i), .Z(w20o));
	IVHSP inv040 (.A(w20o), .Z(w21i));
	IVHSP inv041 (.A(w21i), .Z(w21o));
	IVHSP inv042 (.A(w21o), .Z(w22i));
	IVHSP inv043 (.A(w22i), .Z(w22o));
	IVHSP inv044 (.A(w22o), .Z(w23i));
	IVHSP inv045 (.A(w23i), .Z(w23o));
	IVHSP inv046 (.A(w23o), .Z(w24i));
	IVHSP inv047 (.A(w24i), .Z(w24o));
	IVHSP inv048 (.A(w24o), .Z(w25i));
	IVHSP inv049 (.A(w25i), .Z(w25o));
	IVHSP inv050 (.A(w25o), .Z(w26i));
	IVHSP inv051 (.A(w26i), .Z(w26o));
	IVHSP inv052 (.A(w26o), .Z(w27i));
	IVHSP inv053 (.A(w27i), .Z(w27o));
	IVHSP inv054 (.A(w27o), .Z(w28i));
	IVHSP inv055 (.A(w28i), .Z(w28o));
	IVHSP inv056 (.A(w28o), .Z(w29i));
	IVHSP inv057 (.A(w29i), .Z(w29o));
	IVHSP inv058 (.A(w29o), .Z(w30i));
	IVHSP inv059 (.A(w30i), .Z(w30o));
	IVHSP inv060 (.A(w30o), .Z(w31i));
	IVHSP inv061 (.A(w31i), .Z(w31o));
	IVHSP inv062 (.A(w31o), .Z(w32i));
	IVHSP inv063 (.A(w32i), .Z(w32o));
	IVHSP inv064 (.A(w32o), .Z(w33i));
	IVHSP inv065 (.A(w33i), .Z(w33o));
	IVHSP inv066 (.A(w33o), .Z(w34i));
	IVHSP inv067 (.A(w34i), .Z(w34o));
	IVHSP inv068 (.A(w34o), .Z(w35i));
	IVHSP inv069 (.A(w35i), .Z(w35o));
	IVHSP inv070 (.A(w35o), .Z(w36i));
	IVHSP inv071 (.A(w36i), .Z(w36o));
	IVHSP inv072 (.A(w36o), .Z(w37i));
	IVHSP inv073 (.A(w37i), .Z(w37o));
	IVHSP inv074 (.A(w37o), .Z(w38i));
	IVHSP inv075 (.A(w38i), .Z(w38o));
	IVHSP inv076 (.A(w38o), .Z(w39i));
	IVHSP inv077 (.A(w39i), .Z(w39o));
	IVHSP inv078 (.A(w39o), .Z(w40i));
	IVHSP inv079 (.A(w40i), .Z(w40o));
	IVHSP inv080 (.A(w40o), .Z(w41i));
	IVHSP inv081 (.A(w41i), .Z(w41o));
	IVHSP inv082 (.A(w41o), .Z(w42i));
	IVHSP inv083 (.A(w42i), .Z(w42o));
	IVHSP inv084 (.A(w42o), .Z(w43i));
	IVHSP inv085 (.A(w43i), .Z(w43o));
	IVHSP inv086 (.A(w43o), .Z(w44i));
	IVHSP inv087 (.A(w44i), .Z(w44o));
	IVHSP inv088 (.A(w44o), .Z(w45i));
	IVHSP inv089 (.A(w45i), .Z(w45o));
	IVHSP inv090 (.A(w45o), .Z(w46i));
	IVHSP inv091 (.A(w46i), .Z(w46o));
	IVHSP inv092 (.A(w46o), .Z(w47i));
	IVHSP inv093 (.A(w47i), .Z(w47o));
	IVHSP inv094 (.A(w47o), .Z(w48i));
	IVHSP inv095 (.A(w48i), .Z(w48o));
	IVHSP inv096 (.A(w48o), .Z(w49i));
	IVHSP inv097 (.A(w49i), .Z(w49o));
	IVHSP inv098 (.A(w49o), .Z(w50i));
	IVHSP inv099 (.A(w50i), .Z(w50o));
	IVHSP inv100 (.A(w50o), .Z(w51i));
	IVHSP inv101 (.A(w51i), .Z(w51o));
	IVHSP inv102 (.A(w51o), .Z(w52i));
	IVHSP inv103 (.A(w52i), .Z(w52o));
	IVHSP inv104 (.A(w52o), .Z(w53i));
	IVHSP inv105 (.A(w53i), .Z(w53o));
	IVHSP inv106 (.A(w53o), .Z(wo));

	ND2HSP nand0 (.A(wo), .B(rst_n), .Z(wi));
	FD2HSP ff0 (.D(diff_lb), .CP(wo), .Q(clk_out), .QN(diff_lb), .CD(rst_n));

endmodule
